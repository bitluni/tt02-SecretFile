module secretFile (
    input [7:0] io_in,
    output reg [7:0] io_out
);

wire clk = io_in[0];

reg [9:0] index;

always@(posedge clk) begin
	if(index == 10'd816)
		index <= 10'd0;
	else
		index <= index + 1'd1;
	case(index)
		10'b0000000000: io_out <= 8'b01000111;
		10'b0000000001: io_out <= 8'b01001001;
		10'b0000000010: io_out <= 8'b01000110;
		10'b0000000011: io_out <= 8'b00111000;
		10'b0000000100: io_out <= 8'b00111001;
		10'b0000000101: io_out <= 8'b01100001;
		10'b0000000110: io_out <= 8'b00100000;
		10'b0000001000: io_out <= 8'b00100000;
		10'b0000001010: io_out <= 8'b11110010;
		10'b0000001011: io_out <= 8'b00000101;
		10'b0000001101: io_out <= 8'b00110001;
		10'b0000001110: io_out <= 8'b00101100;
		10'b0000001111: io_out <= 8'b00100000;
		10'b0000010000: io_out <= 8'b01011010;
		10'b0000010001: io_out <= 8'b01001000;
		10'b0000010010: io_out <= 8'b01000001;
		10'b0000010011: io_out <= 8'b10011001;
		10'b0000010100: io_out <= 8'b01101011;
		10'b0000010101: io_out <= 8'b01101001;
		10'b0000010110: io_out <= 8'b10001111;
		10'b0000010111: io_out <= 8'b01111110;
		10'b0000011000: io_out <= 8'b10000100;
		10'b0000011001: io_out <= 8'b10011111;
		10'b0000011010: io_out <= 8'b10011101;
		10'b0000011011: io_out <= 8'b10101101;
		10'b0000011100: io_out <= 8'b10101010;
		10'b0000011101: io_out <= 8'b10110001;
		10'b0000011110: io_out <= 8'b11001111;
		10'b0000011111: io_out <= 8'b10111001;
		10'b0000100000: io_out <= 8'b11000000;
		10'b0000100001: io_out <= 8'b11100000;
		10'b0000100101: io_out <= 8'b00100001;
		10'b0000100110: io_out <= 8'b11111111;
		10'b0000100111: io_out <= 8'b00001011;
		10'b0000101000: io_out <= 8'b01001110;
		10'b0000101001: io_out <= 8'b01000101;
		10'b0000101010: io_out <= 8'b01010100;
		10'b0000101011: io_out <= 8'b01010011;
		10'b0000101100: io_out <= 8'b01000011;
		10'b0000101101: io_out <= 8'b01000001;
		10'b0000101110: io_out <= 8'b01010000;
		10'b0000101111: io_out <= 8'b01000101;
		10'b0000110000: io_out <= 8'b00110010;
		10'b0000110001: io_out <= 8'b00101110;
		10'b0000110010: io_out <= 8'b00110000;
		10'b0000110011: io_out <= 8'b00000011;
		10'b0000110100: io_out <= 8'b00000001;
		10'b0000111000: io_out <= 8'b00100001;
		10'b0000111001: io_out <= 8'b11111001;
		10'b0000111010: io_out <= 8'b00000100;
		10'b0000111011: io_out <= 8'b00000100;
		10'b0000111100: io_out <= 8'b00010110;
		10'b0001000000: io_out <= 8'b00100001;
		10'b0001000001: io_out <= 8'b11111110;
		10'b0001000010: io_out <= 8'b00101001;
		10'b0001000011: io_out <= 8'b01001110;
		10'b0001000100: io_out <= 8'b01100101;
		10'b0001000101: io_out <= 8'b01110110;
		10'b0001000110: io_out <= 8'b01100101;
		10'b0001000111: io_out <= 8'b01110010;
		10'b0001001000: io_out <= 8'b00100000;
		10'b0001001001: io_out <= 8'b01100111;
		10'b0001001010: io_out <= 8'b01101111;
		10'b0001001011: io_out <= 8'b01101110;
		10'b0001001100: io_out <= 8'b01101110;
		10'b0001001101: io_out <= 8'b01100001;
		10'b0001001110: io_out <= 8'b00100000;
		10'b0001001111: io_out <= 8'b01100111;
		10'b0001010000: io_out <= 8'b01101001;
		10'b0001010001: io_out <= 8'b01110110;
		10'b0001010010: io_out <= 8'b01100101;
		10'b0001010011: io_out <= 8'b00100000;
		10'b0001010100: io_out <= 8'b01111001;
		10'b0001010101: io_out <= 8'b01101111;
		10'b0001010110: io_out <= 8'b01110101;
		10'b0001010111: io_out <= 8'b00100000;
		10'b0001011000: io_out <= 8'b01110101;
		10'b0001011001: io_out <= 8'b01110000;
		10'b0001011010: io_out <= 8'b00100001;
		10'b0001011011: io_out <= 8'b00100000;
		10'b0001011100: io_out <= 8'b01100010;
		10'b0001011101: io_out <= 8'b01101001;
		10'b0001011110: io_out <= 8'b01110100;
		10'b0001011111: io_out <= 8'b01101100;
		10'b0001100000: io_out <= 8'b01110101;
		10'b0001100001: io_out <= 8'b01101110;
		10'b0001100010: io_out <= 8'b01101001;
		10'b0001100011: io_out <= 8'b00100000;
		10'b0001100100: io_out <= 8'b01110111;
		10'b0001100101: io_out <= 8'b01100001;
		10'b0001100110: io_out <= 8'b01110011;
		10'b0001100111: io_out <= 8'b00100000;
		10'b0001101000: io_out <= 8'b01101000;
		10'b0001101001: io_out <= 8'b01100101;
		10'b0001101010: io_out <= 8'b01110010;
		10'b0001101011: io_out <= 8'b01100101;
		10'b0001101101: io_out <= 8'b00101100;
		10'b0001110010: io_out <= 8'b00100000;
		10'b0001110100: io_out <= 8'b00100000;
		10'b0001110111: io_out <= 8'b00000011;
		10'b0001111000: io_out <= 8'b10101110;
		10'b0001111001: io_out <= 8'b01011000;
		10'b0001111010: io_out <= 8'b10111010;
		10'b0001111011: io_out <= 8'b10111100;
		10'b0001111100: io_out <= 8'b11110100;
		10'b0001111101: io_out <= 8'b11010000;
		10'b0001111110: io_out <= 8'b11000101;
		10'b0001111111: io_out <= 8'b01101000;
		10'b0010000000: io_out <= 8'b01011010;
		10'b0010000001: io_out <= 8'b10111101;
		10'b0010000010: io_out <= 8'b10010010;
		10'b0010000011: io_out <= 8'b10101010;
		10'b0010000100: io_out <= 8'b01001001;
		10'b0010000101: io_out <= 8'b10110000;
		10'b0010000110: io_out <= 8'b01101111;
		10'b0010000111: io_out <= 8'b01011100;
		10'b0010001000: io_out <= 8'b00010110;
		10'b0010001001: io_out <= 8'b01110110;
		10'b0010001010: io_out <= 8'b00010110;
		10'b0010001011: io_out <= 8'b00111000;
		10'b0010001100: io_out <= 8'b00001001;
		10'b0010001101: io_out <= 8'b11000010;
		10'b0010001110: io_out <= 8'b00011000;
		10'b0010001111: io_out <= 8'b10010110;
		10'b0010010000: io_out <= 8'b10100010;
		10'b0010010001: io_out <= 8'b00010000;
		10'b0010010010: io_out <= 8'b10111100;
		10'b0010010011: io_out <= 8'b10101001;
		10'b0010010100: io_out <= 8'b00111000;
		10'b0010010101: io_out <= 8'b01111101;
		10'b0010010110: io_out <= 8'b10100110;
		10'b0010010111: io_out <= 8'b11111011;
		10'b0010011000: io_out <= 8'b11000010;
		10'b0010011001: io_out <= 8'b11101010;
		10'b0010011010: io_out <= 8'b01000011;
		10'b0010011011: io_out <= 8'b01100011;
		10'b0010011100: io_out <= 8'b00010000;
		10'b0010011101: io_out <= 8'b11101010;
		10'b0010011110: io_out <= 8'b10100011;
		10'b0010011111: io_out <= 8'b10100100;
		10'b0010100000: io_out <= 8'b11001101;
		10'b0010100001: io_out <= 8'b10001010;
		10'b0010100010: io_out <= 8'b11010101;
		10'b0010100011: io_out <= 8'b11111011;
		10'b0010100100: io_out <= 8'b00000001;
		10'b0010100101: io_out <= 8'b01110011;
		10'b0010100110: io_out <= 8'b10101100;
		10'b0010100111: io_out <= 8'b10001100;
		10'b0010101000: io_out <= 8'b11110001;
		10'b0010101001: io_out <= 8'b10001000;
		10'b0010101010: io_out <= 8'b01001100;
		10'b0010101011: io_out <= 8'b00010110;
		10'b0010101100: io_out <= 8'b01111111;
		10'b0010101101: io_out <= 8'b11001000;
		10'b0010101110: io_out <= 8'b00100000;
		10'b0010101111: io_out <= 8'b11110001;
		10'b0010110000: io_out <= 8'b10110001;
		10'b0010110001: io_out <= 8'b11001100;
		10'b0010110010: io_out <= 8'b01101001;
		10'b0010110011: io_out <= 8'b01100110;
		10'b0010110100: io_out <= 8'b01000010;
		10'b0010110101: io_out <= 8'b10000010;
		10'b0010110110: io_out <= 8'b10110001;
		10'b0010110111: io_out <= 8'b00101001;
		10'b0010111000: io_out <= 8'b11001011;
		10'b0010111001: io_out <= 8'b00111110;
		10'b0010111010: io_out <= 8'b01100011;
		10'b0010111011: io_out <= 8'b01010001;
		10'b0010111100: io_out <= 8'b10101111;
		10'b0010111101: io_out <= 8'b10011000;
		10'b0010111110: io_out <= 8'b00010000;
		10'b0010111111: io_out <= 8'b11111000;
		10'b0011000000: io_out <= 8'b10010101;
		10'b0011000001: io_out <= 8'b10100011;
		10'b0011000010: io_out <= 8'b11101000;
		10'b0011000011: io_out <= 8'b10110010;
		10'b0011000100: io_out <= 8'b00101111;
		10'b0011000111: io_out <= 8'b11100000;
		10'b0011001000: io_out <= 8'b10110000;
		10'b0011001001: io_out <= 8'b01010111;
		10'b0011001010: io_out <= 8'b10001110;
		10'b0011001011: io_out <= 8'b01111010;
		10'b0011001100: io_out <= 8'b11100000;
		10'b0011001101: io_out <= 8'b01101010;
		10'b0011001110: io_out <= 8'b11011011;
		10'b0011001111: io_out <= 8'b00000011;
		10'b0011010000: io_out <= 8'b11110000;
		10'b0011010001: io_out <= 8'b10101110;
		10'b0011010010: io_out <= 8'b00101011;
		10'b0011010011: io_out <= 8'b00000101;
		10'b0011010100: io_out <= 8'b01100100;
		10'b0011010101: io_out <= 8'b11011011;
		10'b0011010110: io_out <= 8'b11011011;
		10'b0011010111: io_out <= 8'b01100111;
		10'b0011011000: io_out <= 8'b01101000;
		10'b0011011001: io_out <= 8'b01011010;
		10'b0011011010: io_out <= 8'b01101100;
		10'b0011011011: io_out <= 8'b01111000;
		10'b0011011100: io_out <= 8'b00101000;
		10'b0011011101: io_out <= 8'b00101111;
		10'b0011011110: io_out <= 8'b01111111;
		10'b0011011111: io_out <= 8'b01110111;
		10'b0011100000: io_out <= 8'b10000010;
		10'b0011100001: io_out <= 8'b00110111;
		10'b0011100010: io_out <= 8'b10000000;
		10'b0011100011: io_out <= 8'b10001011;
		10'b0011100100: io_out <= 8'b10001000;
		10'b0011100101: io_out <= 8'b10000000;
		10'b0011100110: io_out <= 8'b01011100;
		10'b0011100111: io_out <= 8'b00000010;
		10'b0011101000: io_out <= 8'b01101110;
		10'b0011101001: io_out <= 8'b01110111;
		10'b0011101010: io_out <= 8'b10001101;
		10'b0011101011: io_out <= 8'b10001110;
		10'b0011101100: io_out <= 8'b01111000;
		10'b0011101101: io_out <= 8'b01010001;
		10'b0011101110: io_out <= 8'b10010001;
		10'b0011101111: io_out <= 8'b01111111;
		10'b0011110000: io_out <= 8'b00110111;
		10'b0011110001: io_out <= 8'b01111110;
		10'b0011110010: io_out <= 8'b10010101;
		10'b0011110011: io_out <= 8'b10000010;
		10'b0011110100: io_out <= 8'b10001000;
		10'b0011110101: io_out <= 8'b10010100;
		10'b0011110110: io_out <= 8'b10011100;
		10'b0011110111: io_out <= 8'b01101000;
		10'b0011111000: io_out <= 8'b10011110;
		10'b0011111001: io_out <= 8'b10000111;
		10'b0011111010: io_out <= 8'b10001110;
		10'b0011111011: io_out <= 8'b01110110;
		10'b0011111100: io_out <= 8'b00000011;
		10'b0011111101: io_out <= 8'b01101001;
		10'b0011111110: io_out <= 8'b10011001;
		10'b0011111111: io_out <= 8'b10100011;
		10'b0100000000: io_out <= 8'b10100100;
		10'b0100000001: io_out <= 8'b01101110;
		10'b0100000010: io_out <= 8'b10100111;
		10'b0100000011: io_out <= 8'b10010011;
		10'b0100000100: io_out <= 8'b10011011;
		10'b0100000101: io_out <= 8'b10100100;
		10'b0100000110: io_out <= 8'b10010110;
		10'b0100000111: io_out <= 8'b01010110;
		10'b0100001000: io_out <= 8'b10101110;
		10'b0100001001: io_out <= 8'b10011111;
		10'b0100001010: io_out <= 8'b10100000;
		10'b0100001011: io_out <= 8'b10110001;
		10'b0100001100: io_out <= 8'b10101000;
		10'b0100001101: io_out <= 8'b10101110;
		10'b0100001110: io_out <= 8'b10110100;
		10'b0100001111: io_out <= 8'b00101010;
		10'b0100010000: io_out <= 8'b01110101;
		10'b0100010001: io_out <= 8'b10101000;
		10'b0100010010: io_out <= 8'b10101010;
		10'b0100010011: io_out <= 8'b10001111;
		10'b0100010100: io_out <= 8'b00111001;
		10'b0100010101: io_out <= 8'b01101011;
		10'b0100010110: io_out <= 8'b10111100;
		10'b0100010111: io_out <= 8'b10101111;
		10'b0100011000: io_out <= 8'b01010110;
		10'b0100011001: io_out <= 8'b00111110;
		10'b0100011010: io_out <= 8'b11000000;
		10'b0100011011: io_out <= 8'b11000001;
		10'b0100011100: io_out <= 8'b11000010;
		10'b0100011101: io_out <= 8'b10011000;
		10'b0100011110: io_out <= 8'b10001100;
		10'b0100011111: io_out <= 8'b11000100;
		10'b0100100000: io_out <= 8'b10100110;
		10'b0100100001: io_out <= 8'b10110101;
		10'b0100100010: io_out <= 8'b10110110;
		10'b0100100011: io_out <= 8'b10110111;
		10'b0100100100: io_out <= 8'b10001001;
		10'b0100100101: io_out <= 8'b00001111;
		10'b0100100110: io_out <= 8'b00001001;
		10'b0100101000: io_out <= 8'b00100001;
		10'b0100101001: io_out <= 8'b11111001;
		10'b0100101010: io_out <= 8'b00000100;
		10'b0100101011: io_out <= 8'b00000101;
		10'b0100101100: io_out <= 8'b00010110;
		10'b0100110000: io_out <= 8'b00101100;
		10'b0100110101: io_out <= 8'b00100000;
		10'b0100110111: io_out <= 8'b00100000;
		10'b0100111001: io_out <= 8'b10000010;
		10'b0100111010: io_out <= 8'b10101010;
		10'b0100111011: io_out <= 8'b10110001;
		10'b0100111100: io_out <= 8'b11001111;
		10'b0100111101: io_out <= 8'b00110001;
		10'b0100111110: io_out <= 8'b00101011;
		10'b0100111111: io_out <= 8'b00011101;
		10'b0101000000: io_out <= 8'b01011001;
		10'b0101000001: io_out <= 8'b01000110;
		10'b0101000010: io_out <= 8'b00111110;
		10'b0101000011: io_out <= 8'b10011000;
		10'b0101000100: io_out <= 8'b01101010;
		10'b0101000101: io_out <= 8'b01100110;
		10'b0101000110: io_out <= 8'b10000111;
		10'b0101000111: io_out <= 8'b01111100;
		10'b0101001000: io_out <= 8'b10000010;
		10'b0101001001: io_out <= 8'b10011110;
		10'b0101001010: io_out <= 8'b10011001;
		10'b0101001011: io_out <= 8'b10101001;
		10'b0101001100: io_out <= 8'b10101010;
		10'b0101001101: io_out <= 8'b10110010;
		10'b0101001110: io_out <= 8'b11010000;
		10'b0101010010: io_out <= 8'b00000011;
		10'b0101010011: io_out <= 8'b11100101;
		10'b0101010100: io_out <= 8'b01101000;
		10'b0101010101: io_out <= 8'b10111010;
		10'b0101010110: io_out <= 8'b01101100;
		10'b0101010111: io_out <= 8'b11110101;
		10'b0101011000: io_out <= 8'b00110000;
		10'b0101011001: io_out <= 8'b11001010;
		10'b0101011010: io_out <= 8'b00000010;
		10'b0101011011: io_out <= 8'b01000000;
		10'b0101011100: io_out <= 8'b10101011;
		10'b0101011101: io_out <= 8'b11001101;
		10'b0101011110: io_out <= 8'b11010100;
		10'b0101011111: io_out <= 8'b11111101;
		10'b0101100000: io_out <= 8'b10000110;
		10'b0101100001: io_out <= 8'b10011111;
		10'b0101100010: io_out <= 8'b10010100;
		10'b0101100011: io_out <= 8'b10100101;
		10'b0101100100: io_out <= 8'b01101101;
		10'b0101100101: io_out <= 8'b01100010;
		10'b0101100110: io_out <= 8'b00100011;
		10'b0101100111: io_out <= 8'b00001101;
		10'b0101101000: io_out <= 8'b01000010;
		10'b0101101001: io_out <= 8'b00101010;
		10'b0101101010: io_out <= 8'b00001100;
		10'b0101101011: io_out <= 8'b10100000;
		10'b0101101100: io_out <= 8'b10000010;
		10'b0101101101: io_out <= 8'b10111001;
		10'b0101101110: io_out <= 8'b10100010;
		10'b0101101111: io_out <= 8'b01111000;
		10'b0101110000: io_out <= 8'b10101010;
		10'b0101110001: io_out <= 8'b00101011;
		10'b0101110010: io_out <= 8'b11111000;
		10'b0101110011: io_out <= 8'b10001100;
		10'b0101110100: io_out <= 8'b11001011;
		10'b0101110101: io_out <= 8'b11000110;
		10'b0101110110: io_out <= 8'b00010100;
		10'b0101110111: io_out <= 8'b10001110;
		10'b0101111000: io_out <= 8'b11100111;
		10'b0101111001: io_out <= 8'b01111111;
		10'b0101111010: io_out <= 8'b00110110;
		10'b0101111011: io_out <= 8'b11010010;
		10'b0101111100: io_out <= 8'b11001011;
		10'b0101111101: io_out <= 8'b11010100;
		10'b0101111110: io_out <= 8'b11111011;
		10'b0101111111: io_out <= 8'b00000001;
		10'b0110000000: io_out <= 8'b00100101;
		10'b0110000001: io_out <= 8'b10010101;
		10'b0110000010: io_out <= 8'b00010000;
		10'b0110000011: io_out <= 8'b00101100;
		10'b0110000100: io_out <= 8'b10100011;
		10'b0110000101: io_out <= 8'b00101000;
		10'b0110000110: io_out <= 8'b00011000;
		10'b0110000111: io_out <= 8'b00111111;
		10'b0110001000: io_out <= 8'b10001110;
		10'b0110001001: io_out <= 8'b00010110;
		10'b0110001010: io_out <= 8'b10101110;
		10'b0110001011: io_out <= 8'b01100100;
		10'b0110001100: io_out <= 8'b01111010;
		10'b0110001101: io_out <= 8'b10110110;
		10'b0110001110: io_out <= 8'b00100000;
		10'b0110001111: io_out <= 8'b00010111;
		10'b0110010000: io_out <= 8'b00010011;
		10'b0110010001: io_out <= 8'b11000100;
		10'b0110010010: io_out <= 8'b00111010;
		10'b0110010011: io_out <= 8'b01110001;
		10'b0110010100: io_out <= 8'b10001100;
		10'b0110010101: io_out <= 8'b10101000;
		10'b0110010110: io_out <= 8'b01011010;
		10'b0110010111: io_out <= 8'b10011110;
		10'b0110011000: io_out <= 8'b11010011;
		10'b0110011001: io_out <= 8'b01100111;
		10'b0110011010: io_out <= 8'b11100011;
		10'b0110011011: io_out <= 8'b01111001;
		10'b0110011100: io_out <= 8'b10011001;
		10'b0110011101: io_out <= 8'b00001011;
		10'b0110011110: io_out <= 8'b01110011;
		10'b0110011111: io_out <= 8'b10000111;
		10'b0110100000: io_out <= 8'b01101100;
		10'b0110100001: io_out <= 8'b10001011;
		10'b0110100010: io_out <= 8'b00110010;
		10'b0110100011: io_out <= 8'b10000100;
		10'b0110100100: io_out <= 8'b11101110;
		10'b0110100101: io_out <= 8'b11101000;
		10'b0110100110: io_out <= 8'b10101111;
		10'b0110100111: io_out <= 8'b01111100;
		10'b0110101000: io_out <= 8'b11011011;
		10'b0110101001: io_out <= 8'b01100001;
		10'b0110101010: io_out <= 8'b10100011;
		10'b0110101011: io_out <= 8'b11100011;
		10'b0110101100: io_out <= 8'b11110001;
		10'b0110101101: io_out <= 8'b10111100;
		10'b0110101110: io_out <= 8'b00001100;
		10'b0110101111: io_out <= 8'b10010111;
		10'b0110110000: io_out <= 8'b11010000;
		10'b0110110001: io_out <= 8'b01010000;
		10'b0110110010: io_out <= 8'b00111110;
		10'b0110110011: io_out <= 8'b00110100;
		10'b0110110100: io_out <= 8'b00100000;
		10'b0110110101: io_out <= 8'b01110000;
		10'b0110110110: io_out <= 8'b01111000;
		10'b0110110111: io_out <= 8'b00110100;
		10'b0110111000: io_out <= 8'b00000001;
		10'b0110111001: io_out <= 8'b00101011;
		10'b0110111010: io_out <= 8'b00101011;
		10'b0110111011: io_out <= 8'b00101100;
		10'b0110111100: io_out <= 8'b00101001;
		10'b0110111101: io_out <= 8'b00000001;
		10'b0110111110: io_out <= 8'b10000111;
		10'b0110111111: io_out <= 8'b00110101;
		10'b0111000000: io_out <= 8'b00010000;
		10'b0111000001: io_out <= 8'b10000100;
		10'b0111000010: io_out <= 8'b00111100;
		10'b0111000011: io_out <= 8'b00000100;
		10'b0111000100: io_out <= 8'b10001101;
		10'b0111000101: io_out <= 8'b00000010;
		10'b0111000110: io_out <= 8'b10010011;
		10'b0111000111: io_out <= 8'b00000010;
		10'b0111001000: io_out <= 8'b00001111;
		10'b0111001001: io_out <= 8'b10010100;
		10'b0111001010: io_out <= 8'b10001100;
		10'b0111001011: io_out <= 8'b10001100;
		10'b0111001100: io_out <= 8'b10001110;
		10'b0111001101: io_out <= 8'b00001111;
		10'b0111001110: io_out <= 8'b00011100;
		10'b0111001111: io_out <= 8'b10000101;
		10'b0111010000: io_out <= 8'b10010100;
		10'b0111010001: io_out <= 8'b10001011;
		10'b0111010010: io_out <= 8'b10011010;
		10'b0111010011: io_out <= 8'b00101001;
		10'b0111010100: io_out <= 8'b00101000;
		10'b0111010101: io_out <= 8'b10011001;
		10'b0111010110: io_out <= 8'b10011001;
		10'b0111010111: io_out <= 8'b10010110;
		10'b0111011000: io_out <= 8'b10001111;
		10'b0111011010: io_out <= 8'b00010011;
		10'b0111011011: io_out <= 8'b10100000;
		10'b0111011100: io_out <= 8'b10100101;
		10'b0111011101: io_out <= 8'b00101000;
		10'b0111011110: io_out <= 8'b10101010;
		10'b0111011111: io_out <= 8'b10100001;
		10'b0111100000: io_out <= 8'b10100110;
		10'b0111100001: io_out <= 8'b00010001;
		10'b0111100010: io_out <= 8'b00011100;
		10'b0111100011: io_out <= 8'b10010111;
		10'b0111100100: io_out <= 8'b10100100;
		10'b0111100101: io_out <= 8'b10101110;
		10'b0111100110: io_out <= 8'b10101101;
		10'b0111100111: io_out <= 8'b10010011;
		10'b0111101000: io_out <= 8'b01110100;
		10'b0111101001: io_out <= 8'b01001110;
		10'b0111101010: io_out <= 8'b10110011;
		10'b0111101011: io_out <= 8'b10110100;
		10'b0111101100: io_out <= 8'b10111001;
		10'b0111101101: io_out <= 8'b10001001;
		10'b0111101110: io_out <= 8'b01101101;
		10'b0111101111: io_out <= 8'b10110010;
		10'b0111110000: io_out <= 8'b10111001;
		10'b0111110001: io_out <= 8'b10010011;
		10'b0111110010: io_out <= 8'b10111001;
		10'b0111110011: io_out <= 8'b01101100;
		10'b0111110100: io_out <= 8'b01011101;
		10'b0111110101: io_out <= 8'b10111110;
		10'b0111110110: io_out <= 8'b10100101;
		10'b0111110111: io_out <= 8'b00110100;
		10'b0111111000: io_out <= 8'b10011000;
		10'b0111111001: io_out <= 8'b10101011;
		10'b0111111010: io_out <= 8'b01000111;
		10'b0111111011: io_out <= 8'b00100000;
		10'b0111111100: io_out <= 8'b10101101;
		10'b0111111101: io_out <= 8'b10001001;
		10'b0111111110: io_out <= 8'b00101010;
		10'b0111111111: io_out <= 8'b10111111;
		10'b1000000000: io_out <= 8'b10001000;
		10'b1000000001: io_out <= 8'b00010011;
		10'b1000000010: io_out <= 8'b00011100;
		10'b1000000011: io_out <= 8'b11001101;
		10'b1000000100: io_out <= 8'b10000111;
		10'b1000000101: io_out <= 8'b00011110;
		10'b1000000110: io_out <= 8'b10011111;
		10'b1000000111: io_out <= 8'b10110101;
		10'b1000001000: io_out <= 8'b10010011;
		10'b1000001001: io_out <= 8'b00101100;
		10'b1000001010: io_out <= 8'b00110110;
		10'b1000001011: io_out <= 8'b10101010;
		10'b1000001100: io_out <= 8'b11001100;
		10'b1000001101: io_out <= 8'b10001101;
		10'b1000001110: io_out <= 8'b10111111;
		10'b1000001111: io_out <= 8'b10101011;
		10'b1000010000: io_out <= 8'b10100111;
		10'b1000010001: io_out <= 8'b01001001;
		10'b1000010010: io_out <= 8'b11000111;
		10'b1000010011: io_out <= 8'b10111011;
		10'b1000010100: io_out <= 8'b11100001;
		10'b1000010101: io_out <= 8'b11001110;
		10'b1000010110: io_out <= 8'b11011111;
		10'b1000010111: io_out <= 8'b10101000;
		10'b1000011000: io_out <= 8'b00000101;
		10'b1000011001: io_out <= 8'b10000110;
		10'b1000011010: io_out <= 8'b10100100;
		10'b1000011011: io_out <= 8'b11010110;
		10'b1000011100: io_out <= 8'b10110011;
		10'b1000011101: io_out <= 8'b11011000;
		10'b1000011110: io_out <= 8'b11100101;
		10'b1000011111: io_out <= 8'b00011101;
		10'b1000100000: io_out <= 8'b11100011;
		10'b1000100001: io_out <= 8'b11101010;
		10'b1000100010: io_out <= 8'b10100101;
		10'b1000100011: io_out <= 8'b10110111;
		10'b1000100100: io_out <= 8'b11000100;
		10'b1000100101: io_out <= 8'b10100001;
		10'b1000100110: io_out <= 8'b11011101;
		10'b1000100111: io_out <= 8'b10011010;
		10'b1000101000: io_out <= 8'b11110010;
		10'b1000101001: io_out <= 8'b11100111;
		10'b1000101010: io_out <= 8'b10110011;
		10'b1000101011: io_out <= 8'b11100011;
		10'b1000101100: io_out <= 8'b11000101;
		10'b1000101101: io_out <= 8'b11110111;
		10'b1000101110: io_out <= 8'b11110011;
		10'b1000101111: io_out <= 8'b11011100;
		10'b1000110000: io_out <= 8'b10111011;
		10'b1000110001: io_out <= 8'b11101100;
		10'b1000110010: io_out <= 8'b11110010;
		10'b1000110011: io_out <= 8'b11011110;
		10'b1000110100: io_out <= 8'b11101001;
		10'b1000110101: io_out <= 8'b10110011;
		10'b1000110110: io_out <= 8'b00010111;
		10'b1000110111: io_out <= 8'b00100001;
		10'b1000111000: io_out <= 8'b00000001;
		10'b1000111010: io_out <= 8'b00100001;
		10'b1000111011: io_out <= 8'b11111001;
		10'b1000111100: io_out <= 8'b00000100;
		10'b1000111101: io_out <= 8'b00000101;
		10'b1000111110: io_out <= 8'b00010110;
		10'b1001000010: io_out <= 8'b00101100;
		10'b1001000111: io_out <= 8'b00100000;
		10'b1001001001: io_out <= 8'b00100000;
		10'b1001001011: io_out <= 8'b10000010;
		10'b1001001100: io_out <= 8'b00110001;
		10'b1001001101: io_out <= 8'b00101100;
		10'b1001001110: io_out <= 8'b00100000;
		10'b1001001111: io_out <= 8'b00110000;
		10'b1001010000: io_out <= 8'b00101011;
		10'b1001010001: io_out <= 8'b00011111;
		10'b1001010010: io_out <= 8'b01011001;
		10'b1001010011: io_out <= 8'b01001001;
		10'b1001010100: io_out <= 8'b01000010;
		10'b1001010101: io_out <= 8'b10011001;
		10'b1001010110: io_out <= 8'b01101000;
		10'b1001010111: io_out <= 8'b01100101;
		10'b1001011000: io_out <= 8'b10011111;
		10'b1001011001: io_out <= 8'b10011010;
		10'b1001011010: io_out <= 8'b10101001;
		10'b1001011011: io_out <= 8'b10101010;
		10'b1001011100: io_out <= 8'b10110001;
		10'b1001011101: io_out <= 8'b11001111;
		10'b1001011110: io_out <= 8'b10101101;
		10'b1001011111: io_out <= 8'b10110011;
		10'b1001100000: io_out <= 8'b11010000;
		10'b1001100100: io_out <= 8'b00000011;
		10'b1001100101: io_out <= 8'b11001000;
		10'b1001100110: io_out <= 8'b01101000;
		10'b1001100111: io_out <= 8'b10111010;
		10'b1001101000: io_out <= 8'b10101100;
		10'b1001101001: io_out <= 8'b11110100;
		10'b1001101010: io_out <= 8'b10001111;
		10'b1001101011: io_out <= 8'b11000001;
		10'b1001101100: io_out <= 8'b01001001;
		10'b1001101101: io_out <= 8'b01011010;
		10'b1001101110: io_out <= 8'b10110001;
		10'b1001101111: io_out <= 8'b10001110;
		10'b1001110000: io_out <= 8'b00110110;
		10'b1001110001: io_out <= 8'b00011010;
		10'b1001110010: io_out <= 8'b00010101;
		10'b1001110011: io_out <= 8'b11000000;
		10'b1001110100: io_out <= 8'b00001011;
		10'b1001110101: io_out <= 8'b01010111;
		10'b1001110110: io_out <= 8'b10000101;
		10'b1001110111: io_out <= 8'b00011100;
		10'b1001111000: io_out <= 8'b00011000;
		10'b1001111001: io_out <= 8'b10010010;
		10'b1001111010: io_out <= 8'b01010101;
		10'b1001111011: io_out <= 8'b10000111;
		10'b1001111100: io_out <= 8'b01101010;
		10'b1001111101: io_out <= 8'b10011001;
		10'b1001111110: io_out <= 8'b11111010;
		10'b1001111111: io_out <= 8'b00001100;
		10'b1010000000: io_out <= 8'b10000011;
		10'b1010000010: io_out <= 8'b10001111;
		10'b1010000011: io_out <= 8'b10011011;
		10'b1010000100: io_out <= 8'b01101000;
		10'b1010000110: io_out <= 8'b10101010;
		10'b1010000111: io_out <= 8'b00010011;
		10'b1010001000: io_out <= 8'b00001011;
		10'b1010001001: io_out <= 8'b10111100;
		10'b1010001010: io_out <= 8'b00001100;
		10'b1010001011: io_out <= 8'b01001001;
		10'b1010001100: io_out <= 8'b00110110;
		10'b1010001101: io_out <= 8'b11011010;
		10'b1010001110: io_out <= 8'b01100111;
		10'b1010001111: io_out <= 8'b00010001;
		10'b1010010000: io_out <= 8'b10000011;
		10'b1010010001: io_out <= 8'b00010101;
		10'b1010010010: io_out <= 8'b01011001;
		10'b1010010011: io_out <= 8'b00100010;
		10'b1010010100: io_out <= 8'b11011010;
		10'b1010010101: io_out <= 8'b01000101;
		10'b1010010110: io_out <= 8'b01100010;
		10'b1010010111: io_out <= 8'b01101100;
		10'b1010011000: io_out <= 8'b00100110;
		10'b1010011001: io_out <= 8'b01111111;
		10'b1010011010: io_out <= 8'b00111111;
		10'b1010011011: io_out <= 8'b01010011;
		10'b1010011100: io_out <= 8'b11010011;
		10'b1010011101: io_out <= 8'b00011000;
		10'b1010011110: io_out <= 8'b01001001;
		10'b1010011111: io_out <= 8'b01001010;
		10'b1010100000: io_out <= 8'b10000000;
		10'b1010100001: io_out <= 8'b10111010;
		10'b1010100010: io_out <= 8'b11101001;
		10'b1010100011: io_out <= 8'b10100000;
		10'b1010100100: io_out <= 8'b10000100;
		10'b1010100101: io_out <= 8'b10110100;
		10'b1010100110: io_out <= 8'b10100100;
		10'b1010100111: io_out <= 8'b00001000;
		10'b1010101000: io_out <= 8'b11011010;
		10'b1010101001: io_out <= 8'b00001110;
		10'b1010101010: io_out <= 8'b01110100;
		10'b1010101011: io_out <= 8'b01100010;
		10'b1010101100: io_out <= 8'b11001000;
		10'b1010101101: io_out <= 8'b10010101;
		10'b1010101110: io_out <= 8'b00101001;
		10'b1010101111: io_out <= 8'b01010011;
		10'b1010110000: io_out <= 8'b10101110;
		10'b1010110001: io_out <= 8'b01101101;
		10'b1010110010: io_out <= 8'b00110101;
		10'b1010110011: io_out <= 8'b11010001;
		10'b1010110100: io_out <= 8'b01101110;
		10'b1010110101: io_out <= 8'b11000111;
		10'b1010110110: io_out <= 8'b01000001;
		10'b1010110111: io_out <= 8'b11111000;
		10'b1010111000: io_out <= 8'b10101011;
		10'b1010111001: io_out <= 8'b11101001;
		10'b1010111010: io_out <= 8'b01111011;
		10'b1010111011: io_out <= 8'b00111110;
		10'b1010111100: io_out <= 8'b11001111;
		10'b1010111101: io_out <= 8'b01110011;
		10'b1010111110: io_out <= 8'b01111010;
		10'b1010111111: io_out <= 8'b11001111;
		10'b1011000000: io_out <= 8'b11001110;
		10'b1011000001: io_out <= 8'b11100111;
		10'b1011000010: io_out <= 8'b01101001;
		10'b1011000011: io_out <= 8'b01111001;
		10'b1011000100: io_out <= 8'b00000001;
		10'b1011000101: io_out <= 8'b01111011;
		10'b1011000110: io_out <= 8'b01111100;
		10'b1011000111: io_out <= 8'b00010011;
		10'b1011001000: io_out <= 8'b10000000;
		10'b1011001001: io_out <= 8'b10000001;
		10'b1011001010: io_out <= 8'b01010100;
		10'b1011001011: io_out <= 8'b00000100;
		10'b1011001100: io_out <= 8'b00000010;
		10'b1011001101: io_out <= 8'b00000001;
		10'b1011001110: io_out <= 8'b10001010;
		10'b1011001111: io_out <= 8'b10000110;
		10'b1011010000: io_out <= 8'b10000011;
		10'b1011010001: io_out <= 8'b01100000;
		10'b1011010010: io_out <= 8'b10001001;
		10'b1011010011: io_out <= 8'b10001011;
		10'b1011010100: io_out <= 8'b00000010;
		10'b1011010101: io_out <= 8'b01100000;
		10'b1011010110: io_out <= 8'b01101111;
		10'b1011010111: io_out <= 8'b10001111;
		10'b1011011000: io_out <= 8'b10010000;
		10'b1011011001: io_out <= 8'b10001101;
		10'b1011011010: io_out <= 8'b10010100;
		10'b1011011011: io_out <= 8'b10001010;
		10'b1011011100: io_out <= 8'b00111101;
		10'b1011011101: io_out <= 8'b10011001;
		10'b1011011110: io_out <= 8'b10001011;
		10'b1011011111: io_out <= 8'b10011000;
		10'b1011100000: io_out <= 8'b10000011;
		10'b1011100001: io_out <= 8'b00000011;
		10'b1011100010: io_out <= 8'b10011011;
		10'b1011100011: io_out <= 8'b10010000;
		10'b1011100100: io_out <= 8'b10011001;
		10'b1011100101: io_out <= 8'b10010111;
		10'b1011100110: io_out <= 8'b10000001;
		10'b1011100111: io_out <= 8'b10000011;
		10'b1011101000: io_out <= 8'b10100010;
		10'b1011101001: io_out <= 8'b10100000;
		10'b1011101010: io_out <= 8'b10000101;
		10'b1011101011: io_out <= 8'b10011011;
		10'b1011101100: io_out <= 8'b10010001;
		10'b1011101101: io_out <= 8'b00011010;
		10'b1011101110: io_out <= 8'b00010100;
		10'b1011101111: io_out <= 8'b10100101;
		10'b1011110000: io_out <= 8'b10011000;
		10'b1011110001: io_out <= 8'b10011010;
		10'b1011110010: io_out <= 8'b10011111;
		10'b1011110011: io_out <= 8'b01101111;
		10'b1011110100: io_out <= 8'b01001111;
		10'b1011110101: io_out <= 8'b10101100;
		10'b1011110110: io_out <= 8'b10000001;
		10'b1011110111: io_out <= 8'b10100001;
		10'b1011111000: io_out <= 8'b10100111;
		10'b1011111001: io_out <= 8'b10101001;
		10'b1011111010: io_out <= 8'b10110001;
		10'b1011111011: io_out <= 8'b10011111;
		10'b1011111100: io_out <= 8'b10101000;
		10'b1011111101: io_out <= 8'b00111101;
		10'b1011111110: io_out <= 8'b01000110;
		10'b1011111111: io_out <= 8'b10001111;
		10'b1100000000: io_out <= 8'b10110110;
		10'b1100000001: io_out <= 8'b01001001;
		10'b1100000010: io_out <= 8'b10110010;
		10'b1100000011: io_out <= 8'b10110011;
		10'b1100000100: io_out <= 8'b01111110;
		10'b1100000101: io_out <= 8'b00110000;
		10'b1100000110: io_out <= 8'b10111100;
		10'b1100000111: io_out <= 8'b01111101;
		10'b1100001000: io_out <= 8'b10111000;
		10'b1100001001: io_out <= 8'b10100110;
		10'b1100001010: io_out <= 8'b11000001;
		10'b1100001011: io_out <= 8'b10010100;
		10'b1100001100: io_out <= 8'b10110000;
		10'b1100001101: io_out <= 8'b00100010;
		10'b1100001110: io_out <= 8'b10111111;
		10'b1100001111: io_out <= 8'b10110011;
		10'b1100010000: io_out <= 8'b10101101;
		10'b1100010001: io_out <= 8'b11000011;
		10'b1100010010: io_out <= 8'b01110110;
		10'b1100010011: io_out <= 8'b10100111;
		10'b1100010100: io_out <= 8'b10111000;
		10'b1100010101: io_out <= 8'b11010000;
		10'b1100010110: io_out <= 8'b10011000;
		10'b1100010111: io_out <= 8'b11001001;
		10'b1100011000: io_out <= 8'b00100010;
		10'b1100011001: io_out <= 8'b10111011;
		10'b1100011010: io_out <= 8'b11000101;
		10'b1100011011: io_out <= 8'b11010010;
		10'b1100011100: io_out <= 8'b00111100;
		10'b1100011101: io_out <= 8'b10011101;
		10'b1100011110: io_out <= 8'b11000010;
		10'b1100011111: io_out <= 8'b11010111;
		10'b1100100000: io_out <= 8'b10010100;
		10'b1100100001: io_out <= 8'b01110101;
		10'b1100100010: io_out <= 8'b11011010;
		10'b1100100011: io_out <= 8'b00110001;
		10'b1100100100: io_out <= 8'b11000101;
		10'b1100100101: io_out <= 8'b10000001;
		10'b1100100110: io_out <= 8'b10010101;
		10'b1100100111: io_out <= 8'b10001101;
		10'b1100101000: io_out <= 8'b10010010;
		10'b1100101001: io_out <= 8'b11100000;
		10'b1100101010: io_out <= 8'b11010001;
		10'b1100101011: io_out <= 8'b10100111;
		10'b1100101100: io_out <= 8'b01111100;
		10'b1100101101: io_out <= 8'b00001001;
		10'b1100101111: io_out <= 8'b00111011;
		default: io_out <= 8'b00000000;
	endcase;
end

endmodule
