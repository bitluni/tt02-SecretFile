module option23 (
    input [7:0] io_in,
    output reg [7:0] io_out
);

parameter WORD_COUNT = 20;

wire clk = io_in[0];
wire [6:0] din = io_in[7:1];

reg [2:0] counter;
reg [7 * WORD_COUNT - 1: 0] buffer;

always@(posedge clk) begin
    if(din == 7'b1111111) begin
        if(!buffer[6]) begin
            io_out <= {1'b0, buffer[5:0], 1'b0};
            buffer <= {buffer[6: 0], buffer[7 * WORD_COUNT - 1: 7]};
            counter <= 3'd0;
        end else begin
            if(counter == 3'b111) begin
                buffer <= {buffer[6: 0], buffer[7 * WORD_COUNT - 1: 7]};
                counter <= 3'd0;
            end else begin
                counter <= counter + 1'd1;
            end
            case({buffer[5:0], counter[2:0]})
                10'b0010000001: io_out <= 8'b00111110;
                10'b0010000010: io_out <= 8'b01100001;
                10'b0010000011: io_out <= 8'b01010001;
                10'b0010000100: io_out <= 8'b01001001;
                10'b0010000101: io_out <= 8'b01000101;
                10'b0010000110: io_out <= 8'b00111110;
                10'b0010001001: io_out <= 8'b01000100;
                10'b0010001010: io_out <= 8'b01000010;
                10'b0010001011: io_out <= 8'b01111111;
                10'b0010001100: io_out <= 8'b01000000;
                10'b0010001101: io_out <= 8'b01000000;
                10'b0010010001: io_out <= 8'b01100010;
                10'b0010010010: io_out <= 8'b01010001;
                10'b0010010011: io_out <= 8'b01010001;
                10'b0010010100: io_out <= 8'b01001001;
                10'b0010010101: io_out <= 8'b01001001;
                10'b0010010110: io_out <= 8'b01100110;
                10'b0010011001: io_out <= 8'b00100010;
                10'b0010011010: io_out <= 8'b01000001;
                10'b0010011011: io_out <= 8'b01001001;
                10'b0010011100: io_out <= 8'b01001001;
                10'b0010011101: io_out <= 8'b01001001;
                10'b0010011110: io_out <= 8'b00110110;
                10'b0010100000: io_out <= 8'b00010000;
                10'b0010100001: io_out <= 8'b00011000;
                10'b0010100010: io_out <= 8'b00010100;
                10'b0010100011: io_out <= 8'b01010010;
                10'b0010100100: io_out <= 8'b01111111;
                10'b0010100101: io_out <= 8'b01010000;
                10'b0010100110: io_out <= 8'b00010000;
                10'b0010101001: io_out <= 8'b00100111;
                10'b0010101010: io_out <= 8'b01000101;
                10'b0010101011: io_out <= 8'b01000101;
                10'b0010101100: io_out <= 8'b01000101;
                10'b0010101101: io_out <= 8'b01000101;
                10'b0010101110: io_out <= 8'b00111001;
                10'b0010110001: io_out <= 8'b00111100;
                10'b0010110010: io_out <= 8'b01001010;
                10'b0010110011: io_out <= 8'b01001001;
                10'b0010110100: io_out <= 8'b01001001;
                10'b0010110101: io_out <= 8'b01001001;
                10'b0010110110: io_out <= 8'b00110000;
                10'b0010111001: io_out <= 8'b00000011;
                10'b0010111010: io_out <= 8'b00000001;
                10'b0010111011: io_out <= 8'b01110001;
                10'b0010111100: io_out <= 8'b00001001;
                10'b0010111101: io_out <= 8'b00000101;
                10'b0010111110: io_out <= 8'b00000011;
                10'b0011000001: io_out <= 8'b00110110;
                10'b0011000010: io_out <= 8'b01001001;
                10'b0011000011: io_out <= 8'b01001001;
                10'b0011000100: io_out <= 8'b01001001;
                10'b0011000101: io_out <= 8'b01001001;
                10'b0011000110: io_out <= 8'b00110110;
                10'b0011001001: io_out <= 8'b00000110;
                10'b0011001010: io_out <= 8'b01001001;
                10'b0011001011: io_out <= 8'b01001001;
                10'b0011001100: io_out <= 8'b01001001;
                10'b0011001101: io_out <= 8'b00101001;
                10'b0011001110: io_out <= 8'b00011110;
                10'b0100001001: io_out <= 8'b01111100;
                10'b0100001010: io_out <= 8'b00010010;
                10'b0100001011: io_out <= 8'b00010001;
                10'b0100001100: io_out <= 8'b00010001;
                10'b0100001101: io_out <= 8'b00010010;
                10'b0100001110: io_out <= 8'b01111100;
                10'b0100010001: io_out <= 8'b01000001;
                10'b0100010010: io_out <= 8'b01111111;
                10'b0100010011: io_out <= 8'b01001001;
                10'b0100010100: io_out <= 8'b01001001;
                10'b0100010101: io_out <= 8'b01001001;
                10'b0100010110: io_out <= 8'b00110110;
                10'b0100011001: io_out <= 8'b00011100;
                10'b0100011010: io_out <= 8'b00100010;
                10'b0100011011: io_out <= 8'b01000001;
                10'b0100011100: io_out <= 8'b01000001;
                10'b0100011101: io_out <= 8'b01000001;
                10'b0100011110: io_out <= 8'b00100010;
                10'b0100100001: io_out <= 8'b01000001;
                10'b0100100010: io_out <= 8'b01111111;
                10'b0100100011: io_out <= 8'b01000001;
                10'b0100100100: io_out <= 8'b01000001;
                10'b0100100101: io_out <= 8'b00100010;
                10'b0100100110: io_out <= 8'b00011100;
                10'b0100101001: io_out <= 8'b01000001;
                10'b0100101010: io_out <= 8'b01111111;
                10'b0100101011: io_out <= 8'b01001001;
                10'b0100101100: io_out <= 8'b01011101;
                10'b0100101101: io_out <= 8'b01000001;
                10'b0100101110: io_out <= 8'b01100011;
                10'b0100110001: io_out <= 8'b01000001;
                10'b0100110010: io_out <= 8'b01111111;
                10'b0100110011: io_out <= 8'b01001001;
                10'b0100110100: io_out <= 8'b00011101;
                10'b0100110101: io_out <= 8'b00000001;
                10'b0100110110: io_out <= 8'b00000011;
                10'b0100111001: io_out <= 8'b00011100;
                10'b0100111010: io_out <= 8'b00100010;
                10'b0100111011: io_out <= 8'b01000001;
                10'b0100111100: io_out <= 8'b01010001;
                10'b0100111101: io_out <= 8'b01010001;
                10'b0100111110: io_out <= 8'b01110010;
                10'b0101000001: io_out <= 8'b01111111;
                10'b0101000010: io_out <= 8'b00001000;
                10'b0101000011: io_out <= 8'b00001000;
                10'b0101000100: io_out <= 8'b00001000;
                10'b0101000101: io_out <= 8'b00001000;
                10'b0101000110: io_out <= 8'b01111111;
                10'b0101001010: io_out <= 8'b01000001;
                10'b0101001011: io_out <= 8'b01111111;
                10'b0101001100: io_out <= 8'b01000001;
                10'b0101010001: io_out <= 8'b00110000;
                10'b0101010010: io_out <= 8'b01000000;
                10'b0101010011: io_out <= 8'b01000000;
                10'b0101010100: io_out <= 8'b01000001;
                10'b0101010101: io_out <= 8'b00111111;
                10'b0101010110: io_out <= 8'b00000001;
                10'b0101011001: io_out <= 8'b01000001;
                10'b0101011010: io_out <= 8'b01111111;
                10'b0101011011: io_out <= 8'b00001000;
                10'b0101011100: io_out <= 8'b00010100;
                10'b0101011101: io_out <= 8'b00100010;
                10'b0101011110: io_out <= 8'b01000001;
                10'b0101011111: io_out <= 8'b01000000;
                10'b0101100001: io_out <= 8'b01000001;
                10'b0101100010: io_out <= 8'b01111111;
                10'b0101100011: io_out <= 8'b01000001;
                10'b0101100100: io_out <= 8'b01000000;
                10'b0101100101: io_out <= 8'b01000000;
                10'b0101100110: io_out <= 8'b01100000;
                10'b0101101001: io_out <= 8'b01111111;
                10'b0101101010: io_out <= 8'b00000001;
                10'b0101101011: io_out <= 8'b00000010;
                10'b0101101100: io_out <= 8'b00000100;
                10'b0101101101: io_out <= 8'b00000010;
                10'b0101101110: io_out <= 8'b00000001;
                10'b0101101111: io_out <= 8'b01111111;
                10'b0101110001: io_out <= 8'b01111111;
                10'b0101110010: io_out <= 8'b00000001;
                10'b0101110011: io_out <= 8'b00000010;
                10'b0101110100: io_out <= 8'b00000100;
                10'b0101110101: io_out <= 8'b00001000;
                10'b0101110110: io_out <= 8'b01111111;
                10'b0101111001: io_out <= 8'b00011100;
                10'b0101111010: io_out <= 8'b00100010;
                10'b0101111011: io_out <= 8'b01000001;
                10'b0101111100: io_out <= 8'b01000001;
                10'b0101111101: io_out <= 8'b00100010;
                10'b0101111110: io_out <= 8'b00011100;
                10'b0110000001: io_out <= 8'b01000001;
                10'b0110000010: io_out <= 8'b01111111;
                10'b0110000011: io_out <= 8'b01001001;
                10'b0110000100: io_out <= 8'b00001001;
                10'b0110000101: io_out <= 8'b00001001;
                10'b0110000110: io_out <= 8'b00000110;
                10'b0110001001: io_out <= 8'b00011110;
                10'b0110001010: io_out <= 8'b00100001;
                10'b0110001011: io_out <= 8'b00100001;
                10'b0110001100: io_out <= 8'b00110001;
                10'b0110001101: io_out <= 8'b00100001;
                10'b0110001110: io_out <= 8'b01011110;
                10'b0110001111: io_out <= 8'b01000000;
                10'b0110010001: io_out <= 8'b01000001;
                10'b0110010010: io_out <= 8'b01111111;
                10'b0110010011: io_out <= 8'b01001001;
                10'b0110010100: io_out <= 8'b00011001;
                10'b0110010101: io_out <= 8'b00101001;
                10'b0110010110: io_out <= 8'b01000110;
                10'b0110011001: io_out <= 8'b00100110;
                10'b0110011010: io_out <= 8'b01001001;
                10'b0110011011: io_out <= 8'b01001001;
                10'b0110011100: io_out <= 8'b01001001;
                10'b0110011101: io_out <= 8'b01001001;
                10'b0110011110: io_out <= 8'b00110010;
                10'b0110100001: io_out <= 8'b00000011;
                10'b0110100010: io_out <= 8'b00000001;
                10'b0110100011: io_out <= 8'b01000001;
                10'b0110100100: io_out <= 8'b01111111;
                10'b0110100101: io_out <= 8'b01000001;
                10'b0110100110: io_out <= 8'b00000001;
                10'b0110100111: io_out <= 8'b00000011;
                10'b0110101001: io_out <= 8'b00111111;
                10'b0110101010: io_out <= 8'b01000000;
                10'b0110101011: io_out <= 8'b01000000;
                10'b0110101100: io_out <= 8'b01000000;
                10'b0110101101: io_out <= 8'b01000000;
                10'b0110101110: io_out <= 8'b00111111;
                10'b0110110001: io_out <= 8'b00001111;
                10'b0110110010: io_out <= 8'b00010000;
                10'b0110110011: io_out <= 8'b00100000;
                10'b0110110100: io_out <= 8'b01000000;
                10'b0110110101: io_out <= 8'b00100000;
                10'b0110110110: io_out <= 8'b00010000;
                10'b0110110111: io_out <= 8'b00001111;
                10'b0110111001: io_out <= 8'b00111111;
                10'b0110111010: io_out <= 8'b01000000;
                10'b0110111011: io_out <= 8'b01000000;
                10'b0110111100: io_out <= 8'b00111000;
                10'b0110111101: io_out <= 8'b01000000;
                10'b0110111110: io_out <= 8'b01000000;
                10'b0110111111: io_out <= 8'b00111111;
                10'b0111000001: io_out <= 8'b01000001;
                10'b0111000010: io_out <= 8'b00100010;
                10'b0111000011: io_out <= 8'b00010100;
                10'b0111000100: io_out <= 8'b00001000;
                10'b0111000101: io_out <= 8'b00010100;
                10'b0111000110: io_out <= 8'b00100010;
                10'b0111000111: io_out <= 8'b01000001;
                10'b0111001001: io_out <= 8'b00000001;
                10'b0111001010: io_out <= 8'b00000010;
                10'b0111001011: io_out <= 8'b01000100;
                10'b0111001100: io_out <= 8'b01111000;
                10'b0111001101: io_out <= 8'b01000100;
                10'b0111001110: io_out <= 8'b00000010;
                10'b0111001111: io_out <= 8'b00000001;
                10'b0111010001: io_out <= 8'b01000011;
                10'b0111010010: io_out <= 8'b01100001;
                10'b0111010011: io_out <= 8'b01010001;
                10'b0111010100: io_out <= 8'b01001001;
                10'b0111010101: io_out <= 8'b01000101;
                10'b0111010110: io_out <= 8'b01000011;
                10'b0111010111: io_out <= 8'b01100001;
                default: io_out <= 8'b00000000;
            endcase;
        end
    end else begin
        buffer <= {din, buffer[7 * WORD_COUNT - 1: 7]};
        io_out <= 8'd0;
        counter <= 3'd0;
    end
end

endmodule
