module charRom (
    input [5:0] face,
    input [2:0] index,
    output [7:0] col
);

assign col = rom[{face,index}];

localparam [511:0][7:0] rom = {
8'b10000000,
8'b10000000,
8'b10000000,
8'b10000000,
8'b10000000,
8'b10000000,
8'b10000000,
8'b10000000,
8'b00000000,
8'b00001000,
8'b00000100,
8'b00000010,
8'b00000001,
8'b00000010,
8'b00000100,
8'b00001000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111111,
8'b01000001,
8'b01000001,
8'b01000001,
8'b00000000,
8'b00000000,
8'b01000000,
8'b00100000,
8'b00010000,
8'b00001000,
8'b00000100,
8'b00000010,
8'b00000001,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01000001,
8'b01000001,
8'b01000001,
8'b01111111,
8'b00000000,
8'b01100001,
8'b01000011,
8'b01000101,
8'b01001001,
8'b01010001,
8'b01100001,
8'b01000011,
8'b00000000,
8'b00000001,
8'b00000010,
8'b01000100,
8'b01111000,
8'b01000100,
8'b00000010,
8'b00000001,
8'b00000000,
8'b01000001,
8'b00100010,
8'b00010100,
8'b00001000,
8'b00010100,
8'b00100010,
8'b01000001,
8'b00000000,
8'b00111111,
8'b01000000,
8'b01000000,
8'b00111000,
8'b01000000,
8'b01000000,
8'b00111111,
8'b00000000,
8'b00001111,
8'b00010000,
8'b00100000,
8'b01000000,
8'b00100000,
8'b00010000,
8'b00001111,
8'b00000000,
8'b00000000,
8'b00111111,
8'b01000000,
8'b01000000,
8'b01000000,
8'b01000000,
8'b00111111,
8'b00000000,
8'b00000011,
8'b00000001,
8'b01000001,
8'b01111111,
8'b01000001,
8'b00000001,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00110010,
8'b01001001,
8'b01001001,
8'b01001001,
8'b01001001,
8'b00100110,
8'b00000000,
8'b00000000,
8'b01000110,
8'b00101001,
8'b00011001,
8'b01001001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b01000000,
8'b01011110,
8'b00100001,
8'b00110001,
8'b00100001,
8'b00100001,
8'b00011110,
8'b00000000,
8'b00000000,
8'b00000110,
8'b00001001,
8'b00001001,
8'b01001001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00011100,
8'b00100010,
8'b01000001,
8'b01000001,
8'b00100010,
8'b00011100,
8'b00000000,
8'b00000000,
8'b01111111,
8'b00001000,
8'b00000100,
8'b00000010,
8'b00000001,
8'b01111111,
8'b00000000,
8'b01111111,
8'b00000001,
8'b00000010,
8'b00000100,
8'b00000010,
8'b00000001,
8'b01111111,
8'b00000000,
8'b00000000,
8'b01100000,
8'b01000000,
8'b01000000,
8'b01000001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b01000000,
8'b01000001,
8'b00100010,
8'b00010100,
8'b00001000,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00000001,
8'b00111111,
8'b01000001,
8'b01000000,
8'b01000000,
8'b00110000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01000001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01111111,
8'b00001000,
8'b00001000,
8'b00001000,
8'b00001000,
8'b01111111,
8'b00000000,
8'b00000000,
8'b01110010,
8'b01010001,
8'b01010001,
8'b01000001,
8'b00100010,
8'b00011100,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000001,
8'b00011101,
8'b01001001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b01100011,
8'b01000001,
8'b01011101,
8'b01001001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00011100,
8'b00100010,
8'b01000001,
8'b01000001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00100010,
8'b01000001,
8'b01000001,
8'b01000001,
8'b00100010,
8'b00011100,
8'b00000000,
8'b00000000,
8'b00110110,
8'b01001001,
8'b01001001,
8'b01001001,
8'b01111111,
8'b01000001,
8'b00000000,
8'b00000000,
8'b01111100,
8'b00010010,
8'b00010001,
8'b00010001,
8'b00010010,
8'b01111100,
8'b00000000,
8'b00000000,
8'b00011110,
8'b01010101,
8'b01010101,
8'b01011101,
8'b01000001,
8'b00111110,
8'b00000000,
8'b00000000,
8'b00000110,
8'b00001001,
8'b01010001,
8'b00000001,
8'b00000001,
8'b00000010,
8'b00000000,
8'b00000000,
8'b00001000,
8'b00010100,
8'b00100010,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00100100,
8'b00100100,
8'b00100100,
8'b00100100,
8'b00100100,
8'b00100100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01000001,
8'b00100010,
8'b00010100,
8'b00001000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01100110,
8'b10000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01100110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00011110,
8'b00101001,
8'b01001001,
8'b01001001,
8'b01001001,
8'b00000110,
8'b00000000,
8'b00000000,
8'b00110110,
8'b01001001,
8'b01001001,
8'b01001001,
8'b01001001,
8'b00110110,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000101,
8'b00001001,
8'b01110001,
8'b00000001,
8'b00000011,
8'b00000000,
8'b00000000,
8'b00110000,
8'b01001001,
8'b01001001,
8'b01001001,
8'b01001010,
8'b00111100,
8'b00000000,
8'b00000000,
8'b00111001,
8'b01000101,
8'b01000101,
8'b01000101,
8'b01000101,
8'b00100111,
8'b00000000,
8'b00000000,
8'b00010000,
8'b01010000,
8'b01111111,
8'b01010010,
8'b00010100,
8'b00011000,
8'b00010000,
8'b00000000,
8'b00110110,
8'b01001001,
8'b01001001,
8'b01001001,
8'b01000001,
8'b00100010,
8'b00000000,
8'b00000000,
8'b01100110,
8'b01001001,
8'b01001001,
8'b01010001,
8'b01010001,
8'b01100010,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01000000,
8'b01000000,
8'b01111111,
8'b01000010,
8'b01000100,
8'b00000000,
8'b00000000,
8'b00111110,
8'b01000101,
8'b01001001,
8'b01010001,
8'b01100001,
8'b00111110,
8'b00000000,
8'b00000000,
8'b00000010,
8'b00000100,
8'b00001000,
8'b00010000,
8'b00100000,
8'b01000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01100000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00001000,
8'b00001000,
8'b00001000,
8'b00001000,
8'b00001000,
8'b00001000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01100000,
8'b10000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00001000,
8'b00001000,
8'b00111110,
8'b00001000,
8'b00001000,
8'b00000000,
8'b00000000,
8'b00001000,
8'b00101010,
8'b00011100,
8'b00011100,
8'b00011100,
8'b00101010,
8'b00001000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00011100,
8'b00100010,
8'b01000001,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01000001,
8'b00100010,
8'b00011100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000011,
8'b00000100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b01001000,
8'b01001000,
8'b00110010,
8'b01001101,
8'b01000101,
8'b01001010,
8'b00110000,
8'b00000000,
8'b01100010,
8'b01100100,
8'b00001000,
8'b00010000,
8'b00100110,
8'b01000110,
8'b00000000,
8'b00000000,
8'b00010010,
8'b00101010,
8'b01101011,
8'b01101011,
8'b00101010,
8'b00100100,
8'b00000000,
8'b00000000,
8'b00010100,
8'b01111111,
8'b00010100,
8'b00010100,
8'b01111111,
8'b00010100,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000111,
8'b00000000,
8'b00000000,
8'b00000111,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000110,
8'b01011111,
8'b00000110,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000,
8'b00000000
};

endmodule
