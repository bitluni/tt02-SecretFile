module secretFile (
    input [7:0] io_in,
    output reg [7:0] io_out
);

wire clk = io_in[0];

reg [11:0] index;

always@(posedge clk) begin
	if(index == 11'd2845)
		index <= 0;
	else
		index <= index + 1'd1;
	case(index)
		12'b000000000000: io_out <= 8'b01000111;
		12'b000000000001: io_out <= 8'b01001001;
		12'b000000000010: io_out <= 8'b01000110;
		12'b000000000011: io_out <= 8'b00111000;
		12'b000000000100: io_out <= 8'b00111001;
		12'b000000000101: io_out <= 8'b01100001;
		12'b000000000110: io_out <= 8'b00100000;
		12'b000000001000: io_out <= 8'b00100000;
		12'b000000001010: io_out <= 8'b11110010;
		12'b000000001101: io_out <= 8'b00110001;
		12'b000000001110: io_out <= 8'b00101100;
		12'b000000001111: io_out <= 8'b00100000;
		12'b000000010000: io_out <= 8'b01011010;
		12'b000000010001: io_out <= 8'b01001000;
		12'b000000010010: io_out <= 8'b01000001;
		12'b000000010011: io_out <= 8'b10011001;
		12'b000000010100: io_out <= 8'b01101011;
		12'b000000010101: io_out <= 8'b01101001;
		12'b000000010110: io_out <= 8'b10011111;
		12'b000000010111: io_out <= 8'b10011101;
		12'b000000011000: io_out <= 8'b10101101;
		12'b000000011001: io_out <= 8'b10101010;
		12'b000000011010: io_out <= 8'b10110001;
		12'b000000011011: io_out <= 8'b11001111;
		12'b000000011100: io_out <= 8'b10111001;
		12'b000000011101: io_out <= 8'b11000000;
		12'b000000011110: io_out <= 8'b11100000;
		12'b000000011111: io_out <= 8'b10001111;
		12'b000000100000: io_out <= 8'b01111110;
		12'b000000100001: io_out <= 8'b10000100;
		12'b000000100101: io_out <= 8'b00100001;
		12'b000000100110: io_out <= 8'b11111111;
		12'b000000100111: io_out <= 8'b00001011;
		12'b000000101000: io_out <= 8'b01001110;
		12'b000000101001: io_out <= 8'b01000101;
		12'b000000101010: io_out <= 8'b01010100;
		12'b000000101011: io_out <= 8'b01010011;
		12'b000000101100: io_out <= 8'b01000011;
		12'b000000101101: io_out <= 8'b01000001;
		12'b000000101110: io_out <= 8'b01010000;
		12'b000000101111: io_out <= 8'b01000101;
		12'b000000110000: io_out <= 8'b00110010;
		12'b000000110001: io_out <= 8'b00101110;
		12'b000000110010: io_out <= 8'b00110000;
		12'b000000110011: io_out <= 8'b00000011;
		12'b000000110100: io_out <= 8'b00000001;
		12'b000000111000: io_out <= 8'b00100001;
		12'b000000111001: io_out <= 8'b11111001;
		12'b000000111010: io_out <= 8'b00000100;
		12'b000000111011: io_out <= 8'b00000100;
		12'b000000111100: io_out <= 8'b00001101;
		12'b000001000000: io_out <= 8'b00100001;
		12'b000001000001: io_out <= 8'b11111110;
		12'b000001000010: io_out <= 8'b00101001;
		12'b000001000011: io_out <= 8'b01001110;
		12'b000001000100: io_out <= 8'b01100101;
		12'b000001000101: io_out <= 8'b01110110;
		12'b000001000110: io_out <= 8'b01100101;
		12'b000001000111: io_out <= 8'b01110010;
		12'b000001001000: io_out <= 8'b00100000;
		12'b000001001001: io_out <= 8'b01100111;
		12'b000001001010: io_out <= 8'b01101111;
		12'b000001001011: io_out <= 8'b01101110;
		12'b000001001100: io_out <= 8'b01101110;
		12'b000001001101: io_out <= 8'b01100001;
		12'b000001001110: io_out <= 8'b00100000;
		12'b000001001111: io_out <= 8'b01100111;
		12'b000001010000: io_out <= 8'b01101001;
		12'b000001010001: io_out <= 8'b01110110;
		12'b000001010010: io_out <= 8'b01100101;
		12'b000001010011: io_out <= 8'b00100000;
		12'b000001010100: io_out <= 8'b01111001;
		12'b000001010101: io_out <= 8'b01101111;
		12'b000001010110: io_out <= 8'b01110101;
		12'b000001010111: io_out <= 8'b00100000;
		12'b000001011000: io_out <= 8'b01110101;
		12'b000001011001: io_out <= 8'b01110000;
		12'b000001011010: io_out <= 8'b00100001;
		12'b000001011011: io_out <= 8'b00100000;
		12'b000001011100: io_out <= 8'b01100010;
		12'b000001011101: io_out <= 8'b01101001;
		12'b000001011110: io_out <= 8'b01110100;
		12'b000001011111: io_out <= 8'b01101100;
		12'b000001100000: io_out <= 8'b01110101;
		12'b000001100001: io_out <= 8'b01101110;
		12'b000001100010: io_out <= 8'b01101001;
		12'b000001100011: io_out <= 8'b00100000;
		12'b000001100100: io_out <= 8'b01110111;
		12'b000001100101: io_out <= 8'b01100001;
		12'b000001100110: io_out <= 8'b01110011;
		12'b000001100111: io_out <= 8'b00100000;
		12'b000001101000: io_out <= 8'b01101000;
		12'b000001101001: io_out <= 8'b01100101;
		12'b000001101010: io_out <= 8'b01110010;
		12'b000001101011: io_out <= 8'b01100101;
		12'b000001101101: io_out <= 8'b00101100;
		12'b000001110010: io_out <= 8'b00100000;
		12'b000001110100: io_out <= 8'b00100000;
		12'b000001110111: io_out <= 8'b00000011;
		12'b000001111000: io_out <= 8'b11010100;
		12'b000001111001: io_out <= 8'b01001000;
		12'b000001111010: io_out <= 8'b01010100;
		12'b000001111011: io_out <= 8'b11011010;
		12'b000001111100: io_out <= 8'b11000101;
		12'b000001111101: io_out <= 8'b00100011;
		12'b000001111110: io_out <= 8'b11001010;
		12'b000001111111: io_out <= 8'b01000110;
		12'b000010000000: io_out <= 8'b10100100;
		12'b000010000001: io_out <= 8'b00011101;
		12'b000010000010: io_out <= 8'b10001010;
		12'b000010000011: io_out <= 8'b10101101;
		12'b000010000100: io_out <= 8'b11111100;
		12'b000010000101: io_out <= 8'b11110100;
		12'b000010000110: io_out <= 8'b11000101;
		12'b000010000111: io_out <= 8'b11001101;
		12'b000010001000: io_out <= 8'b00000111;
		12'b000010001001: io_out <= 8'b01110110;
		12'b000010001010: io_out <= 8'b10010100;
		12'b000010001011: io_out <= 8'b00010110;
		12'b000010001100: io_out <= 8'b01111110;
		12'b000010001101: io_out <= 8'b10001010;
		12'b000010001110: io_out <= 8'b00011000;
		12'b000010001111: io_out <= 8'b01110001;
		12'b000010010000: io_out <= 8'b10001110;
		12'b000010010001: io_out <= 8'b10011001;
		12'b000010010010: io_out <= 8'b01011010;
		12'b000010010011: io_out <= 8'b10000010;
		12'b000010010100: io_out <= 8'b00110000;
		12'b000010010101: io_out <= 8'b01010101;
		12'b000010010110: io_out <= 8'b11100010;
		12'b000010010111: io_out <= 8'b11100010;
		12'b000010011000: io_out <= 8'b01101110;
		12'b000010011001: io_out <= 8'b01101111;
		12'b000010011010: io_out <= 8'b00100101;
		12'b000010011011: io_out <= 8'b00000100;
		12'b000010011100: io_out <= 8'b10111100;
		12'b000010011101: io_out <= 8'b01111100;
		12'b000010011110: io_out <= 8'b01111110;
		12'b000010011111: io_out <= 8'b00001111;
		12'b000010100000: io_out <= 8'b00001010;
		12'b000010100001: io_out <= 8'b10001110;
		12'b000010100010: io_out <= 8'b00110110;
		12'b000010100011: io_out <= 8'b11011000;
		12'b000010100100: io_out <= 8'b11110001;
		12'b000010100101: io_out <= 8'b01111010;
		12'b000010100110: io_out <= 8'b00100000;
		12'b000010100111: io_out <= 8'b01010101;
		12'b000010101000: io_out <= 8'b00110000;
		12'b000010101001: io_out <= 8'b11100011;
		12'b000010101010: io_out <= 8'b00100000;
		12'b000010101011: io_out <= 8'b11000110;
		12'b000010101100: io_out <= 8'b10011110;
		12'b000010101101: io_out <= 8'b10110001;
		12'b000010101110: io_out <= 8'b10100100;
		12'b000010101111: io_out <= 8'b01001000;
		12'b000010110000: io_out <= 8'b01100011;
		12'b000010110001: io_out <= 8'b01100010;
		12'b000010110010: io_out <= 8'b01000000;
		12'b000010110011: io_out <= 8'b00100010;
		12'b000010110100: io_out <= 8'b11010000;
		12'b000010110101: io_out <= 8'b01100111;
		12'b000010110110: io_out <= 8'b01101101;
		12'b000010110111: io_out <= 8'b00100110;
		12'b000010111000: io_out <= 8'b10110100;
		12'b000010111001: io_out <= 8'b00111010;
		12'b000010111010: io_out <= 8'b10110011;
		12'b000010111011: io_out <= 8'b00110010;
		12'b000010111100: io_out <= 8'b00010100;
		12'b000010111101: io_out <= 8'b00000110;
		12'b000010111110: io_out <= 8'b11010100;
		12'b000010111111: io_out <= 8'b11011101;
		12'b000011000000: io_out <= 8'b01001000;
		12'b000011000001: io_out <= 8'b11000000;
		12'b000011000010: io_out <= 8'b10101010;
		12'b000011000011: io_out <= 8'b11100100;
		12'b000011000100: io_out <= 8'b11100110;
		12'b000011000101: io_out <= 8'b10010110;
		12'b000011000110: io_out <= 8'b11010010;
		12'b000011000111: io_out <= 8'b01100101;
		12'b000011001000: io_out <= 8'b11010011;
		12'b000011001001: io_out <= 8'b00110100;
		12'b000011001010: io_out <= 8'b11001010;
		12'b000011001011: io_out <= 8'b01011000;
		12'b000011001100: io_out <= 8'b01111010;
		12'b000011001101: io_out <= 8'b10000110;
		12'b000011001110: io_out <= 8'b10100110;
		12'b000011001111: io_out <= 8'b01010111;
		12'b000011010000: io_out <= 8'b11110010;
		12'b000011010001: io_out <= 8'b11011001;
		12'b000011010010: io_out <= 8'b11000111;
		12'b000011010011: io_out <= 8'b01111110;
		12'b000011010100: io_out <= 8'b10011111;
		12'b000011010101: io_out <= 8'b10101111;
		12'b000011010110: io_out <= 8'b00100110;
		12'b000011010111: io_out <= 8'b00011111;
		12'b000011011000: io_out <= 8'b00000001;
		12'b000011011001: io_out <= 8'b01010000;
		12'b000011011010: io_out <= 8'b10000010;
		12'b000011011011: io_out <= 8'b01111101;
		12'b000011011100: io_out <= 8'b01111000;
		12'b000011011101: io_out <= 8'b01110111;
		12'b000011011110: io_out <= 8'b10000010;
		12'b000011011111: io_out <= 8'b01001111;
		12'b000011100000: io_out <= 8'b00000001;
		12'b000011100011: io_out <= 8'b01001000;
		12'b000011100100: io_out <= 8'b00010110;
		12'b000011100101: io_out <= 8'b00111001;
		12'b000011100110: io_out <= 8'b00010101;
		12'b000011100111: io_out <= 8'b01000100;
		12'b000011101000: io_out <= 8'b00010111;
		12'b000011101001: io_out <= 8'b10001000;
		12'b000011101010: io_out <= 8'b00000110;
		12'b000011101011: io_out <= 8'b00111011;
		12'b000011101100: io_out <= 8'b10001011;
		12'b000011101101: io_out <= 8'b10010110;
		12'b000011101110: io_out <= 8'b00000001;
		12'b000011101111: io_out <= 8'b10001110;
		12'b000011110000: io_out <= 8'b01110001;
		12'b000011110001: io_out <= 8'b01111110;
		12'b000011110010: io_out <= 8'b01100111;
		12'b000011110011: io_out <= 8'b10000100;
		12'b000011110100: io_out <= 8'b01010001;
		12'b000011110101: io_out <= 8'b10001010;
		12'b000011110110: io_out <= 8'b10010110;
		12'b000011110111: io_out <= 8'b10001011;
		12'b000011111000: io_out <= 8'b10000100;
		12'b000011111001: io_out <= 8'b10000101;
		12'b000011111010: io_out <= 8'b01011000;
		12'b000011111011: io_out <= 8'b10001010;
		12'b000011111100: io_out <= 8'b10011000;
		12'b000011111101: io_out <= 8'b00110001;
		12'b000011111110: io_out <= 8'b00111100;
		12'b000011111111: io_out <= 8'b10100000;
		12'b000100000000: io_out <= 8'b10010111;
		12'b000100000001: io_out <= 8'b01110111;
		12'b000100000010: io_out <= 8'b00101111;
		12'b000100000011: io_out <= 8'b01000111;
		12'b000100000100: io_out <= 8'b10100001;
		12'b000100000101: io_out <= 8'b10101101;
		12'b000100000110: io_out <= 8'b10101001;
		12'b000100000111: io_out <= 8'b10100001;
		12'b000100001000: io_out <= 8'b01110000;
		12'b000100001001: io_out <= 8'b00101001;
		12'b000100001010: io_out <= 8'b00000010;
		12'b000100001011: io_out <= 8'b10001100;
		12'b000100001100: io_out <= 8'b10010111;
		12'b000100001101: io_out <= 8'b10101111;
		12'b000100001110: io_out <= 8'b10110000;
		12'b000100001111: io_out <= 8'b10011000;
		12'b000100010000: io_out <= 8'b10110010;
		12'b000100010001: io_out <= 8'b01000101;
		12'b000100010010: io_out <= 8'b10101001;
		12'b000100010011: io_out <= 8'b01000111;
		12'b000100010100: io_out <= 8'b10011111;
		12'b000100010101: io_out <= 8'b10111000;
		12'b000100010110: io_out <= 8'b10101011;
		12'b000100010111: io_out <= 8'b00010101;
		12'b000100011000: io_out <= 8'b00000110;
		12'b000100011001: io_out <= 8'b10111100;
		12'b000100011010: io_out <= 8'b10101000;
		12'b000100011011: io_out <= 8'b10110000;
		12'b000100011100: io_out <= 8'b10110001;
		12'b000100011101: io_out <= 8'b10100011;
		12'b000100011110: io_out <= 8'b11000011;
		12'b000100011111: io_out <= 8'b10111110;
		12'b000100100000: io_out <= 8'b11000101;
		12'b000100100001: io_out <= 8'b00000110;
		12'b000100100010: io_out <= 8'b00101010;
		12'b000100100011: io_out <= 8'b10010001;
		12'b000100100100: io_out <= 8'b11001001;
		12'b000100100101: io_out <= 8'b10110111;
		12'b000100100110: io_out <= 8'b11000101;
		12'b000100100111: io_out <= 8'b10111001;
		12'b000100101000: io_out <= 8'b01111101;
		12'b000100101001: io_out <= 8'b11001110;
		12'b000100101010: io_out <= 8'b11000100;
		12'b000100101011: io_out <= 8'b11000101;
		12'b000100101100: io_out <= 8'b10001100;
		12'b000100101101: io_out <= 8'b10100011;
		12'b000100101110: io_out <= 8'b11010011;
		12'b000100101111: io_out <= 8'b11001001;
		12'b000100110000: io_out <= 8'b10111111;
		12'b000100110001: io_out <= 8'b11001100;
		12'b000100110010: io_out <= 8'b00010010;
		12'b000100110011: io_out <= 8'b11011000;
		12'b000100110100: io_out <= 8'b11010101;
		12'b000100110101: io_out <= 8'b11000110;
		12'b000100110110: io_out <= 8'b01110111;
		12'b000100110111: io_out <= 8'b10010101;
		12'b000100111000: io_out <= 8'b10100000;
		12'b000100111001: io_out <= 8'b11010100;
		12'b000100111010: io_out <= 8'b11010000;
		12'b000100111011: io_out <= 8'b01111101;
		12'b000100111100: io_out <= 8'b10001001;
		12'b000100111101: io_out <= 8'b11011110;
		12'b000100111110: io_out <= 8'b11100100;
		12'b000100111111: io_out <= 8'b11100000;
		12'b000101000000: io_out <= 8'b00110001;
		12'b000101000001: io_out <= 8'b11100111;
		12'b000101000010: io_out <= 8'b11101000;
		12'b000101000011: io_out <= 8'b11101001;
		12'b000101000100: io_out <= 8'b11100010;
		12'b000101000101: io_out <= 8'b11011001;
		12'b000101000110: io_out <= 8'b10110000;
		12'b000101000111: io_out <= 8'b11001011;
		12'b000101001000: io_out <= 8'b11010010;
		12'b000101001001: io_out <= 8'b11011000;
		12'b000101001010: io_out <= 8'b11101111;
		12'b000101001011: io_out <= 8'b11011111;
		12'b000101001100: io_out <= 8'b00001001;
		12'b000101001110: io_out <= 8'b00100001;
		12'b000101001111: io_out <= 8'b11111001;
		12'b000101010000: io_out <= 8'b00000100;
		12'b000101010001: io_out <= 8'b00000101;
		12'b000101010010: io_out <= 8'b00001101;
		12'b000101010110: io_out <= 8'b00101100;
		12'b000101011011: io_out <= 8'b00100000;
		12'b000101011101: io_out <= 8'b00100000;
		12'b000101011111: io_out <= 8'b10000010;
		12'b000101100011: io_out <= 8'b00110010;
		12'b000101100100: io_out <= 8'b00101100;
		12'b000101100101: io_out <= 8'b00100000;
		12'b000101100110: io_out <= 8'b01011000;
		12'b000101100111: io_out <= 8'b01000111;
		12'b000101101000: io_out <= 8'b01000000;
		12'b000101101001: io_out <= 8'b10010111;
		12'b000101101010: io_out <= 8'b01101000;
		12'b000101101011: io_out <= 8'b01100100;
		12'b000101101100: io_out <= 8'b10011111;
		12'b000101101101: io_out <= 8'b10011001;
		12'b000101101110: io_out <= 8'b10101000;
		12'b000101101111: io_out <= 8'b10101101;
		12'b000101110000: io_out <= 8'b10110100;
		12'b000101110001: io_out <= 8'b11010000;
		12'b000101110010: io_out <= 8'b10001110;
		12'b000101110011: io_out <= 8'b01111110;
		12'b000101110100: io_out <= 8'b10000101;
		12'b000101111000: io_out <= 8'b00000011;
		12'b000101111001: io_out <= 8'b11111110;
		12'b000101111010: io_out <= 8'b00001000;
		12'b000101111011: io_out <= 8'b10110101;
		12'b000101111100: io_out <= 8'b10111010;
		12'b000101111101: io_out <= 8'b01001110;
		12'b000101111110: io_out <= 8'b00000100;
		12'b000101111111: io_out <= 8'b01001000;
		12'b000110000000: io_out <= 8'b01000000;
		12'b000110000001: io_out <= 8'b10000110;
		12'b000110000010: io_out <= 8'b00011101;
		12'b000110000011: io_out <= 8'b10010001;
		12'b000110000100: io_out <= 8'b01100110;
		12'b000110000101: io_out <= 8'b10100111;
		12'b000110000110: io_out <= 8'b01100100;
		12'b000110000111: io_out <= 8'b10011001;
		12'b000110001000: io_out <= 8'b00011101;
		12'b000110001001: io_out <= 8'b01001000;
		12'b000110001010: io_out <= 8'b00001101;
		12'b000110001011: io_out <= 8'b01000010;
		12'b000110001100: io_out <= 8'b00101001;
		12'b000110001101: io_out <= 8'b00001100;
		12'b000110001110: io_out <= 8'b01100010;
		12'b000110001111: io_out <= 8'b00100011;
		12'b000110010000: io_out <= 8'b00111010;
		12'b000110010001: io_out <= 8'b00011111;
		12'b000110010010: io_out <= 8'b00110011;
		12'b000110010011: io_out <= 8'b01010101;
		12'b000110010100: io_out <= 8'b01100110;
		12'b000110010101: io_out <= 8'b10001001;
		12'b000110010110: io_out <= 8'b01000001;
		12'b000110010111: io_out <= 8'b10110100;
		12'b000110011000: io_out <= 8'b11011011;
		12'b000110011001: io_out <= 8'b01001110;
		12'b000110011010: io_out <= 8'b01101101;
		12'b000110011011: io_out <= 8'b01010001;
		12'b000110011100: io_out <= 8'b01010111;
		12'b000110011101: io_out <= 8'b11010111;
		12'b000110011110: io_out <= 8'b10010101;
		12'b000110011111: io_out <= 8'b10101101;
		12'b000110100000: io_out <= 8'b10011110;
		12'b000110100001: io_out <= 8'b01010000;
		12'b000110100010: io_out <= 8'b01000011;
		12'b000110100011: io_out <= 8'b01000111;
		12'b000110100100: io_out <= 8'b01011000;
		12'b000110100101: io_out <= 8'b11110000;
		12'b000110100110: io_out <= 8'b01111010;
		12'b000110100111: io_out <= 8'b10011000;
		12'b000110101000: io_out <= 8'b10010100;
		12'b000110101001: io_out <= 8'b10010010;
		12'b000110101010: io_out <= 8'b01100101;
		12'b000110101011: io_out <= 8'b00101100;
		12'b000110101100: io_out <= 8'b11101010;
		12'b000110101101: io_out <= 8'b10010000;
		12'b000110101110: io_out <= 8'b10010110;
		12'b000110101111: io_out <= 8'b11011111;
		12'b000110110000: io_out <= 8'b11110010;
		12'b000110110001: io_out <= 8'b00110011;
		12'b000110110010: io_out <= 8'b00110100;
		12'b000110110011: io_out <= 8'b00111110;
		12'b000110110100: io_out <= 8'b10100000;
		12'b000110110101: io_out <= 8'b01000101;
		12'b000110110110: io_out <= 8'b10010000;
		12'b000110110111: io_out <= 8'b10010100;
		12'b000110111000: io_out <= 8'b10011010;
		12'b000110111001: io_out <= 8'b01100011;
		12'b000110111010: io_out <= 8'b00011010;
		12'b000110111011: io_out <= 8'b10110001;
		12'b000110111100: io_out <= 8'b11000000;
		12'b000110111101: io_out <= 8'b01010100;
		12'b000110111110: io_out <= 8'b11010111;
		12'b000110111111: io_out <= 8'b01001010;
		12'b000111000000: io_out <= 8'b00111011;
		12'b000111000001: io_out <= 8'b11001110;
		12'b000111000010: io_out <= 8'b01010110;
		12'b000111000011: io_out <= 8'b01011001;
		12'b000111000100: io_out <= 8'b10011100;
		12'b000111000101: io_out <= 8'b10000111;
		12'b000111000110: io_out <= 8'b01010101;
		12'b000111000111: io_out <= 8'b00101100;
		12'b000111001000: io_out <= 8'b11110111;
		12'b000111001001: io_out <= 8'b11001010;
		12'b000111001010: io_out <= 8'b00111111;
		12'b000111001011: io_out <= 8'b10101011;
		12'b000111001100: io_out <= 8'b10101101;
		12'b000111001101: io_out <= 8'b11101010;
		12'b000111001110: io_out <= 8'b00100100;
		12'b000111001111: io_out <= 8'b00100010;
		12'b000111010000: io_out <= 8'b00001101;
		12'b000111010001: io_out <= 8'b00101111;
		12'b000111010010: io_out <= 8'b00001000;
		12'b000111010011: io_out <= 8'b10010001;
		12'b000111010100: io_out <= 8'b10000101;
		12'b000111010101: io_out <= 8'b10000110;
		12'b000111010110: io_out <= 8'b10011011;
		12'b000111010111: io_out <= 8'b01001001;
		12'b000111011000: io_out <= 8'b00000010;
		12'b000111011001: io_out <= 8'b01111110;
		12'b000111011010: io_out <= 8'b01110101;
		12'b000111011011: io_out <= 8'b00101110;
		12'b000111011100: io_out <= 8'b00011011;
		12'b000111011101: io_out <= 8'b01101110;
		12'b000111011110: io_out <= 8'b00100111;
		12'b000111011111: io_out <= 8'b00111101;
		12'b000111100000: io_out <= 8'b00100101;
		12'b000111100001: io_out <= 8'b00000001;
		12'b000111100010: io_out <= 8'b00100110;
		12'b000111100011: io_out <= 8'b00111111;
		12'b000111100100: io_out <= 8'b01010010;
		12'b000111100101: io_out <= 8'b01000010;
		12'b000111100110: io_out <= 8'b01110110;
		12'b000111100111: io_out <= 8'b00110001;
		12'b000111101000: io_out <= 8'b10000111;
		12'b000111101001: io_out <= 8'b00000100;
		12'b000111101010: io_out <= 8'b10001001;
		12'b000111101011: io_out <= 8'b00000001;
		12'b000111101100: io_out <= 8'b10010100;
		12'b000111101101: io_out <= 8'b00100101;
		12'b000111101110: io_out <= 8'b01010011;
		12'b000111101111: io_out <= 8'b00111000;
		12'b000111110000: io_out <= 8'b10010010;
		12'b000111110001: io_out <= 8'b10010000;
		12'b000111110010: io_out <= 8'b00100111;
		12'b000111110011: io_out <= 8'b10011001;
		12'b000111110100: io_out <= 8'b10010100;
		12'b000111110101: io_out <= 8'b10011101;
		12'b000111110110: io_out <= 8'b10001010;
		12'b000111110111: io_out <= 8'b10001101;
		12'b000111111000: io_out <= 8'b01010101;
		12'b000111111001: io_out <= 8'b00010010;
		12'b000111111010: io_out <= 8'b10011100;
		12'b000111111011: io_out <= 8'b10001010;
		12'b000111111100: io_out <= 8'b10011010;
		12'b000111111101: io_out <= 8'b10010011;
		12'b000111111110: io_out <= 8'b10010101;
		12'b000111111111: io_out <= 8'b10100000;
		12'b001000000000: io_out <= 8'b00111010;
		12'b001000000001: io_out <= 8'b01000100;
		12'b001000000010: io_out <= 8'b00110000;
		12'b001000000011: io_out <= 8'b10010011;
		12'b001000000100: io_out <= 8'b10010000;
		12'b001000000101: io_out <= 8'b00010111;
		12'b001000000110: io_out <= 8'b00000010;
		12'b001000000111: io_out <= 8'b10011101;
		12'b001000001000: io_out <= 8'b10000001;
		12'b001000001001: io_out <= 8'b10001101;
		12'b001000001010: io_out <= 8'b01010010;
		12'b001000001011: io_out <= 8'b00010101;
		12'b001000001100: io_out <= 8'b10001010;
		12'b001000001101: io_out <= 8'b10110000;
		12'b001000001110: io_out <= 8'b00110001;
		12'b001000001111: io_out <= 8'b10101110;
		12'b001000010000: io_out <= 8'b10110000;
		12'b001000010001: io_out <= 8'b00000110;
		12'b001000010010: io_out <= 8'b10100000;
		12'b001000010011: io_out <= 8'b00010100;
		12'b001000010100: io_out <= 8'b01000110;
		12'b001000010101: io_out <= 8'b00100110;
		12'b001000010110: io_out <= 8'b10110110;
		12'b001000010111: io_out <= 8'b00100110;
		12'b001000011000: io_out <= 8'b10111000;
		12'b001000011001: io_out <= 8'b10011101;
		12'b001000011010: io_out <= 8'b10111010;
		12'b001000011011: io_out <= 8'b10110011;
		12'b001000011100: io_out <= 8'b01110101;
		12'b001000011101: io_out <= 8'b10011001;
		12'b001000011110: io_out <= 8'b10101111;
		12'b001000011111: io_out <= 8'b10010101;
		12'b001000100000: io_out <= 8'b10111110;
		12'b001000100001: io_out <= 8'b10000111;
		12'b001000100010: io_out <= 8'b11000111;
		12'b001000100011: io_out <= 8'b10100111;
		12'b001000100100: io_out <= 8'b01001010;
		12'b001000100101: io_out <= 8'b00001101;
		12'b001000100110: io_out <= 8'b00110000;
		12'b001000100111: io_out <= 8'b10011110;
		12'b001000101000: io_out <= 8'b10100100;
		12'b001000101001: io_out <= 8'b11001000;
		12'b001000101010: io_out <= 8'b10100110;
		12'b001000101011: io_out <= 8'b10011111;
		12'b001000101100: io_out <= 8'b11001101;
		12'b001000101101: io_out <= 8'b01000100;
		12'b001000101110: io_out <= 8'b00000110;
		12'b001000101111: io_out <= 8'b11001011;
		12'b001000110000: io_out <= 8'b11001000;
		12'b001000110001: io_out <= 8'b11010000;
		12'b001000110010: io_out <= 8'b10110101;
		12'b001000110011: io_out <= 8'b10110000;
		12'b001000110100: io_out <= 8'b10111011;
		12'b001000110101: io_out <= 8'b10100010;
		12'b001000110110: io_out <= 8'b00000011;
		12'b001000110111: io_out <= 8'b11010000;
		12'b001000111000: io_out <= 8'b11010011;
		12'b001000111001: io_out <= 8'b10110000;
		12'b001000111010: io_out <= 8'b10011110;
		12'b001000111011: io_out <= 8'b10010110;
		12'b001000111100: io_out <= 8'b01111101;
		12'b001000111101: io_out <= 8'b10100011;
		12'b001000111110: io_out <= 8'b11010010;
		12'b001000111111: io_out <= 8'b11011010;
		12'b001001000000: io_out <= 8'b11011010;
		12'b001001000001: io_out <= 8'b10000001;
		12'b001001000010: io_out <= 8'b00101001;
		12'b001001000011: io_out <= 8'b00110100;
		12'b001001000100: io_out <= 8'b00010110;
		12'b001001000101: io_out <= 8'b11001011;
		12'b001001000110: io_out <= 8'b10111110;
		12'b001001000111: io_out <= 8'b11101000;
		12'b001001001000: io_out <= 8'b10011110;
		12'b001001001001: io_out <= 8'b11011101;
		12'b001001001010: io_out <= 8'b00010100;
		12'b001001001011: io_out <= 8'b00000110;
		12'b001001001100: io_out <= 8'b00010110;
		12'b001001001101: io_out <= 8'b10110110;
		12'b001001001110: io_out <= 8'b11110000;
		12'b001001001111: io_out <= 8'b11100011;
		12'b001001010000: io_out <= 8'b00010000;
		12'b001001010001: io_out <= 8'b01100010;
		12'b001001010010: io_out <= 8'b00010000;
		12'b001001010011: io_out <= 8'b11000001;
		12'b001001010100: io_out <= 8'b11011000;
		12'b001001010101: io_out <= 8'b11110000;
		12'b001001010110: io_out <= 8'b10110001;
		12'b001001010111: io_out <= 8'b11011101;
		12'b001001011000: io_out <= 8'b00111100;
		12'b001001011001: io_out <= 8'b01011000;
		12'b001001011010: io_out <= 8'b11011101;
		12'b001001011011: io_out <= 8'b11111011;
		12'b001001011100: io_out <= 8'b01010100;
		12'b001001011101: io_out <= 8'b01000110;
		12'b001001011110: io_out <= 8'b00001001;
		12'b001001011111: io_out <= 8'b00001101;
		12'b001001100000: io_out <= 8'b00011001;
		12'b001001100001: io_out <= 8'b10101111;
		12'b001001100010: io_out <= 8'b11000010;
		12'b001001100011: io_out <= 8'b11100001;
		12'b001001100100: io_out <= 8'b00010011;
		12'b001001100101: io_out <= 8'b11000100;
		12'b001001100110: io_out <= 8'b11110000;
		12'b001001100111: io_out <= 8'b11011001;
		12'b001001101000: io_out <= 8'b00111011;
		12'b001001101001: io_out <= 8'b01110100;
		12'b001001101010: io_out <= 8'b00001100;
		12'b001001101011: io_out <= 8'b10110101;
		12'b001001101100: io_out <= 8'b10010100;
		12'b001001101101: io_out <= 8'b11010001;
		12'b001001101110: io_out <= 8'b01110100;
		12'b001001101111: io_out <= 8'b11101111;
		12'b001001110000: io_out <= 8'b01011111;
		12'b001001110001: io_out <= 8'b11000011;
		12'b001001110010: io_out <= 8'b10001001;
		12'b001001110011: io_out <= 8'b10010000;
		12'b001001110100: io_out <= 8'b00101010;
		12'b001001110101: io_out <= 8'b11010010;
		12'b001001110110: io_out <= 8'b01001000;
		12'b001001111001: io_out <= 8'b00100001;
		12'b001001111010: io_out <= 8'b11111001;
		12'b001001111011: io_out <= 8'b00000100;
		12'b001001111100: io_out <= 8'b00000101;
		12'b001001111101: io_out <= 8'b00001101;
		12'b001010000001: io_out <= 8'b00101100;
		12'b001010000110: io_out <= 8'b00100000;
		12'b001010001000: io_out <= 8'b00100000;
		12'b001010001010: io_out <= 8'b10000010;
		12'b001010001110: io_out <= 8'b00110001;
		12'b001010001111: io_out <= 8'b00101011;
		12'b001010010000: io_out <= 8'b00011101;
		12'b001010010001: io_out <= 8'b01011001;
		12'b001010010010: io_out <= 8'b01000110;
		12'b001010010011: io_out <= 8'b00111110;
		12'b001010010100: io_out <= 8'b10011000;
		12'b001010010101: io_out <= 8'b01101010;
		12'b001010010110: io_out <= 8'b01100110;
		12'b001010010111: io_out <= 8'b10011100;
		12'b001010011000: io_out <= 8'b10011010;
		12'b001010011001: io_out <= 8'b10101010;
		12'b001010011010: io_out <= 8'b10101010;
		12'b001010011011: io_out <= 8'b10110010;
		12'b001010011100: io_out <= 8'b11010000;
		12'b001010011101: io_out <= 8'b10000111;
		12'b001010011110: io_out <= 8'b01111100;
		12'b001010011111: io_out <= 8'b10000010;
		12'b001010100011: io_out <= 8'b00000011;
		12'b001010100100: io_out <= 8'b11101101;
		12'b001010100101: io_out <= 8'b01011000;
		12'b001010100110: io_out <= 8'b10111010;
		12'b001010100111: io_out <= 8'b00000101;
		12'b001010101000: io_out <= 8'b01011110;
		12'b001010101001: io_out <= 8'b00100100;
		12'b001010101010: io_out <= 8'b11001010;
		12'b001010101011: io_out <= 8'b01001001;
		12'b001010101100: io_out <= 8'b11001001;
		12'b001010101101: io_out <= 8'b01100011;
		12'b001010101110: io_out <= 8'b00010111;
		12'b001010101111: io_out <= 8'b00111011;
		12'b001010110000: io_out <= 8'b00010111;
		12'b001010110001: io_out <= 8'b10000111;
		12'b001010110010: io_out <= 8'b10101111;
		12'b001010110011: io_out <= 8'b00010110;
		12'b001010110100: io_out <= 8'b10100000;
		12'b001010110101: io_out <= 8'b01101100;
		12'b001010110110: io_out <= 8'b00011001;
		12'b001010110111: io_out <= 8'b01000011;
		12'b001010111000: io_out <= 8'b00001101;
		12'b001010111001: io_out <= 8'b01000010;
		12'b001010111010: io_out <= 8'b00101010;
		12'b001010111011: io_out <= 8'b00001100;
		12'b001010111100: io_out <= 8'b11100000;
		12'b001010111101: io_out <= 8'b00101000;
		12'b001010111110: io_out <= 8'b10111010;
		12'b001010111111: io_out <= 8'b00101110;
		12'b001011000000: io_out <= 8'b11011001;
		12'b001011000001: io_out <= 8'b10101001;
		12'b001011000010: io_out <= 8'b00101011;
		12'b001011000011: io_out <= 8'b00011000;
		12'b001011000100: io_out <= 8'b00110101;
		12'b001011000101: io_out <= 8'b00101111;
		12'b001011000110: io_out <= 8'b10011110;
		12'b001011000111: io_out <= 8'b01000011;
		12'b001011001000: io_out <= 8'b10010000;
		12'b001011001001: io_out <= 8'b11100111;
		12'b001011001010: io_out <= 8'b01111111;
		12'b001011001011: io_out <= 8'b00110110;
		12'b001011001100: io_out <= 8'b11010010;
		12'b001011001101: io_out <= 8'b01100101;
		12'b001011001110: io_out <= 8'b01000111;
		12'b001011001111: io_out <= 8'b11101000;
		12'b001011010000: io_out <= 8'b11111101;
		12'b001011010001: io_out <= 8'b10000000;
		12'b001011010010: io_out <= 8'b00010100;
		12'b001011010011: io_out <= 8'b11001110;
		12'b001011010100: io_out <= 8'b01110000;
		12'b001011010101: io_out <= 8'b01100111;
		12'b001011010110: io_out <= 8'b00111010;
		12'b001011010111: io_out <= 8'b01111110;
		12'b001011011000: io_out <= 8'b00100000;
		12'b001011011001: io_out <= 8'b00101101;
		12'b001011011010: io_out <= 8'b10011100;
		12'b001011011011: io_out <= 8'b10101110;
		12'b001011011100: io_out <= 8'b10100001;
		12'b001011011101: io_out <= 8'b00100011;
		12'b001011011110: io_out <= 8'b00111000;
		12'b001011011111: io_out <= 8'b01011011;
		12'b001011100000: io_out <= 8'b00010010;
		12'b001011100001: io_out <= 8'b11000110;
		12'b001011100010: io_out <= 8'b01010100;
		12'b001011100011: io_out <= 8'b00110100;
		12'b001011100100: io_out <= 8'b10111001;
		12'b001011100101: io_out <= 8'b01010110;
		12'b001011100110: io_out <= 8'b01111000;
		12'b001011100111: io_out <= 8'b00011011;
		12'b001011101000: io_out <= 8'b10101101;
		12'b001011101001: io_out <= 8'b11101001;
		12'b001011101010: io_out <= 8'b01100110;
		12'b001011101011: io_out <= 8'b11110101;
		12'b001011101100: io_out <= 8'b11011001;
		12'b001011101101: io_out <= 8'b10001010;
		12'b001011101110: io_out <= 8'b00111100;
		12'b001011101111: io_out <= 8'b10110001;
		12'b001011110000: io_out <= 8'b01001001;
		12'b001011110001: io_out <= 8'b11010001;
		12'b001011110010: io_out <= 8'b00110001;
		12'b001011110011: io_out <= 8'b11011011;
		12'b001011110100: io_out <= 8'b10100000;
		12'b001011110101: io_out <= 8'b10011010;
		12'b001011110110: io_out <= 8'b11110000;
		12'b001011110111: io_out <= 8'b00001101;
		12'b001011111000: io_out <= 8'b11111010;
		12'b001011111001: io_out <= 8'b00111011;
		12'b001011111010: io_out <= 8'b11001111;
		12'b001011111011: io_out <= 8'b00010111;
		12'b001011111100: io_out <= 8'b00010011;
		12'b001011111101: io_out <= 8'b01110110;
		12'b001011111110: io_out <= 8'b10111011;
		12'b001011111111: io_out <= 8'b01011100;
		12'b001100000000: io_out <= 8'b00111111;
		12'b001100000001: io_out <= 8'b00001011;
		12'b001100000010: io_out <= 8'b10100001;
		12'b001100000011: io_out <= 8'b00010010;
		12'b001100000100: io_out <= 8'b00110100;
		12'b001100000101: io_out <= 8'b00101000;
		12'b001100000110: io_out <= 8'b00111110;
		12'b001100000111: io_out <= 8'b00110100;
		12'b001100001000: io_out <= 8'b00100000;
		12'b001100001001: io_out <= 8'b01111111;
		12'b001100001010: io_out <= 8'b10000000;
		12'b001100001011: io_out <= 8'b00110100;
		12'b001100001100: io_out <= 8'b00000001;
		12'b001100001101: io_out <= 8'b00101011;
		12'b001100001110: io_out <= 8'b00101011;
		12'b001100001111: io_out <= 8'b00101100;
		12'b001100010000: io_out <= 8'b00101001;
		12'b001100010001: io_out <= 8'b00000001;
		12'b001100010010: io_out <= 8'b10001010;
		12'b001100010011: io_out <= 8'b00000010;
		12'b001100010100: io_out <= 8'b00000110;
		12'b001100010101: io_out <= 8'b00010011;
		12'b001100010110: io_out <= 8'b10000111;
		12'b001100010111: io_out <= 8'b01000101;
		12'b001100011000: io_out <= 8'b00000110;
		12'b001100011001: io_out <= 8'b10010000;
		12'b001100011010: io_out <= 8'b00000010;
		12'b001100011011: io_out <= 8'b10010111;
		12'b001100011100: io_out <= 8'b00000010;
		12'b001100011101: io_out <= 8'b00010001;
		12'b001100011110: io_out <= 8'b10011000;
		12'b001100011111: io_out <= 8'b10001111;
		12'b001100100000: io_out <= 8'b10001111;
		12'b001100100001: io_out <= 8'b10010001;
		12'b001100100010: io_out <= 8'b10010011;
		12'b001100100011: io_out <= 8'b00011100;
		12'b001100100100: io_out <= 8'b10001000;
		12'b001100100101: io_out <= 8'b10011000;
		12'b001100100110: io_out <= 8'b10001110;
		12'b001100100111: io_out <= 8'b10011110;
		12'b001100101000: io_out <= 8'b00101001;
		12'b001100101001: io_out <= 8'b00101000;
		12'b001100101010: io_out <= 8'b10011101;
		12'b001100101011: io_out <= 8'b10011101;
		12'b001100101100: io_out <= 8'b10011010;
		12'b001100101101: io_out <= 8'b00010010;
		12'b001100101110: io_out <= 8'b00011100;
		12'b001100101111: io_out <= 8'b00010100;
		12'b001100110000: io_out <= 8'b10100100;
		12'b001100110001: io_out <= 8'b10101001;
		12'b001100110010: io_out <= 8'b00101000;
		12'b001100110011: io_out <= 8'b10101110;
		12'b001100110100: io_out <= 8'b10100101;
		12'b001100110101: io_out <= 8'b10101010;
		12'b001100110110: io_out <= 8'b10100000;
		12'b001100111000: io_out <= 8'b10000001;
		12'b001100111001: io_out <= 8'b10101000;
		12'b001100111010: io_out <= 8'b10110010;
		12'b001100111011: io_out <= 8'b10110001;
		12'b001100111100: io_out <= 8'b10010111;
		12'b001100111101: io_out <= 8'b01110110;
		12'b001100111110: io_out <= 8'b00000100;
		12'b001100111111: io_out <= 8'b10010110;
		12'b001101000000: io_out <= 8'b10110111;
		12'b001101000001: io_out <= 8'b10011001;
		12'b001101000010: io_out <= 8'b10111110;
		12'b001101000011: io_out <= 8'b10001100;
		12'b001101000100: io_out <= 8'b01101111;
		12'b001101000101: io_out <= 8'b10011011;
		12'b001101000110: io_out <= 8'b10111110;
		12'b001101000111: io_out <= 8'b10110010;
		12'b001101001000: io_out <= 8'b10111110;
		12'b001101001001: io_out <= 8'b01101110;
		12'b001101001010: io_out <= 8'b01011111;
		12'b001101001011: io_out <= 8'b11000011;
		12'b001101001100: io_out <= 8'b10101000;
		12'b001101001101: io_out <= 8'b00110100;
		12'b001101001110: io_out <= 8'b10111001;
		12'b001101001111: io_out <= 8'b10001100;
		12'b001101010000: io_out <= 8'b00101100;
		12'b001101010001: io_out <= 8'b01100111;
		12'b001101010010: io_out <= 8'b10110001;
		12'b001101010011: io_out <= 8'b10001100;
		12'b001101010100: io_out <= 8'b00101010;
		12'b001101010101: io_out <= 8'b11000100;
		12'b001101010110: io_out <= 8'b10001011;
		12'b001101010111: io_out <= 8'b00010101;
		12'b001101011000: io_out <= 8'b00011011;
		12'b001101011001: io_out <= 8'b00000100;
		12'b001101011010: io_out <= 8'b11010010;
		12'b001101011011: io_out <= 8'b10001010;
		12'b001101011100: io_out <= 8'b00011110;
		12'b001101011101: io_out <= 8'b10100011;
		12'b001101011110: io_out <= 8'b10111001;
		12'b001101011111: io_out <= 8'b10010111;
		12'b001101100000: io_out <= 8'b11001110;
		12'b001101100001: io_out <= 8'b00100000;
		12'b001101100010: io_out <= 8'b10101110;
		12'b001101100011: io_out <= 8'b11010001;
		12'b001101100100: io_out <= 8'b10010000;
		12'b001101100101: io_out <= 8'b11000100;
		12'b001101100110: io_out <= 8'b10101111;
		12'b001101100111: io_out <= 8'b10101011;
		12'b001101101000: io_out <= 8'b11010110;
		12'b001101101001: io_out <= 8'b10011100;
		12'b001101101010: io_out <= 8'b11010011;
		12'b001101101011: io_out <= 8'b11100111;
		12'b001101101100: io_out <= 8'b11100011;
		12'b001101101101: io_out <= 8'b10110011;
		12'b001101101110: io_out <= 8'b00110010;
		12'b001101101111: io_out <= 8'b11010111;
		12'b001101110000: io_out <= 8'b11011000;
		12'b001101110001: io_out <= 8'b10101001;
		12'b001101110010: io_out <= 8'b11101001;
		12'b001101110011: io_out <= 8'b11000100;
		12'b001101110100: io_out <= 8'b11011110;
		12'b001101110101: io_out <= 8'b00010001;
		12'b001101110110: io_out <= 8'b11101100;
		12'b001101110111: io_out <= 8'b10100111;
		12'b001101111000: io_out <= 8'b11001010;
		12'b001101111001: io_out <= 8'b11110000;
		12'b001101111010: io_out <= 8'b10110111;
		12'b001101111011: io_out <= 8'b10110011;
		12'b001101111100: io_out <= 8'b01110110;
		12'b001101111101: io_out <= 8'b11110000;
		12'b001101111110: io_out <= 8'b11011100;
		12'b001101111111: io_out <= 8'b11001010;
		12'b001110000000: io_out <= 8'b01111110;
		12'b001110000001: io_out <= 8'b00011100;
		12'b001110000010: io_out <= 8'b11111011;
		12'b001110000011: io_out <= 8'b11101010;
		12'b001110000100: io_out <= 8'b11110010;
		12'b001110000101: io_out <= 8'b11101101;
		12'b001110000110: io_out <= 8'b11011010;
		12'b001110000111: io_out <= 8'b01110111;
		12'b001110001000: io_out <= 8'b01001111;
		12'b001110001001: io_out <= 8'b10010001;
		12'b001110001010: io_out <= 8'b10100100;
		12'b001110001011: io_out <= 8'b01011101;
		12'b001110001100: io_out <= 8'b10110110;
		12'b001110001101: io_out <= 8'b11101100;
		12'b001110001110: io_out <= 8'b10101001;
		12'b001110001111: io_out <= 8'b10100011;
		12'b001110010000: io_out <= 8'b10010000;
		12'b001110010011: io_out <= 8'b00100001;
		12'b001110010100: io_out <= 8'b11111001;
		12'b001110010101: io_out <= 8'b00000100;
		12'b001110010110: io_out <= 8'b00000101;
		12'b001110010111: io_out <= 8'b00001101;
		12'b001110011011: io_out <= 8'b00101100;
		12'b001110100000: io_out <= 8'b00100000;
		12'b001110100010: io_out <= 8'b00100000;
		12'b001110100100: io_out <= 8'b10000010;
		12'b001110101000: io_out <= 8'b00110001;
		12'b001110101001: io_out <= 8'b00101011;
		12'b001110101010: io_out <= 8'b00011110;
		12'b001110101011: io_out <= 8'b01011100;
		12'b001110101100: io_out <= 8'b01001011;
		12'b001110101101: io_out <= 8'b01000011;
		12'b001110101110: io_out <= 8'b10011001;
		12'b001110101111: io_out <= 8'b01101011;
		12'b001110110000: io_out <= 8'b01101000;
		12'b001110110001: io_out <= 8'b10011111;
		12'b001110110010: io_out <= 8'b10011011;
		12'b001110110011: io_out <= 8'b10101011;
		12'b001110110100: io_out <= 8'b10101101;
		12'b001110110101: io_out <= 8'b10110100;
		12'b001110110110: io_out <= 8'b11010001;
		12'b001110110111: io_out <= 8'b10010101;
		12'b001110111000: io_out <= 8'b01111101;
		12'b001110111001: io_out <= 8'b10000010;
		12'b001110111101: io_out <= 8'b00000011;
		12'b001110111110: io_out <= 8'b11100011;
		12'b001110111111: io_out <= 8'b01011000;
		12'b001111000000: io_out <= 8'b10111010;
		12'b001111000001: io_out <= 8'b00000101;
		12'b001111000010: io_out <= 8'b01011110;
		12'b001111000011: io_out <= 8'b00100100;
		12'b001111000100: io_out <= 8'b11000110;
		12'b001111000101: io_out <= 8'b10100111;
		12'b001111000110: io_out <= 8'b10100100;
		12'b001111000111: io_out <= 8'b10100100;
		12'b001111001000: io_out <= 8'b00001011;
		12'b001111001001: io_out <= 8'b01100111;
		12'b001111001010: io_out <= 8'b11100111;
		12'b001111001011: io_out <= 8'b00100010;
		12'b001111001100: io_out <= 8'b10110011;
		12'b001111001101: io_out <= 8'b00010011;
		12'b001111001110: io_out <= 8'b10100000;
		12'b001111001111: io_out <= 8'b01110000;
		12'b001111010000: io_out <= 8'b11011010;
		12'b001111010001: io_out <= 8'b00000010;
		12'b001111010010: io_out <= 8'b01111010;
		12'b001111010011: io_out <= 8'b11010000;
		12'b001111010100: io_out <= 8'b11101001;
		12'b001111010101: io_out <= 8'b01110001;
		12'b001111010110: io_out <= 8'b11011011;
		12'b001111010111: io_out <= 8'b01001000;
		12'b001111011000: io_out <= 8'b01000110;
		12'b001111011001: io_out <= 8'b11000011;
		12'b001111011010: io_out <= 8'b11100000;
		12'b001111011011: io_out <= 8'b00010001;
		12'b001111011100: io_out <= 8'b10010101;
		12'b001111011101: io_out <= 8'b11011010;
		12'b001111011110: io_out <= 8'b10001000;
		12'b001111011111: io_out <= 8'b00101110;
		12'b001111100000: io_out <= 8'b10011110;
		12'b001111100001: io_out <= 8'b11000110;
		12'b001111100010: io_out <= 8'b10000010;
		12'b001111100011: io_out <= 8'b00010000;
		12'b001111100100: io_out <= 8'b11010011;
		12'b001111100101: io_out <= 8'b10101110;
		12'b001111100110: io_out <= 8'b00010011;
		12'b001111100111: io_out <= 8'b10101001;
		12'b001111101000: io_out <= 8'b10110100;
		12'b001111101001: io_out <= 8'b11101011;
		12'b001111101010: io_out <= 8'b00011001;
		12'b001111101011: io_out <= 8'b00000111;
		12'b001111101100: io_out <= 8'b00011111;
		12'b001111101101: io_out <= 8'b01001011;
		12'b001111101110: io_out <= 8'b10000111;
		12'b001111101111: io_out <= 8'b01010010;
		12'b001111110000: io_out <= 8'b10000010;
		12'b001111110001: io_out <= 8'b11000101;
		12'b001111110010: io_out <= 8'b10011110;
		12'b001111110011: io_out <= 8'b00110010;
		12'b001111110100: io_out <= 8'b10100000;
		12'b001111110101: io_out <= 8'b00001010;
		12'b001111110110: io_out <= 8'b11111000;
		12'b001111110111: io_out <= 8'b00011000;
		12'b001111111000: io_out <= 8'b11101110;
		12'b001111111001: io_out <= 8'b10100000;
		12'b001111111010: io_out <= 8'b00111111;
		12'b001111111011: io_out <= 8'b10011011;
		12'b001111111100: io_out <= 8'b10000100;
		12'b001111111101: io_out <= 8'b01110001;
		12'b001111111110: io_out <= 8'b11010011;
		12'b001111111111: io_out <= 8'b00111001;
		12'b010000000000: io_out <= 8'b10100001;
		12'b010000000001: io_out <= 8'b10000110;
		12'b010000000010: io_out <= 8'b00101001;
		12'b010000000011: io_out <= 8'b10100100;
		12'b010000000100: io_out <= 8'b11001011;
		12'b010000000101: io_out <= 8'b01001101;
		12'b010000000110: io_out <= 8'b01100010;
		12'b010000000111: io_out <= 8'b10100011;
		12'b010000001000: io_out <= 8'b11100010;
		12'b010000001001: io_out <= 8'b01110001;
		12'b010000001010: io_out <= 8'b00111001;
		12'b010000001011: io_out <= 8'b01001001;
		12'b010000001100: io_out <= 8'b11000000;
		12'b010000001101: io_out <= 8'b01001110;
		12'b010000001110: io_out <= 8'b01100111;
		12'b010000001111: io_out <= 8'b11000000;
		12'b010000010000: io_out <= 8'b01011100;
		12'b010000010001: io_out <= 8'b10110101;
		12'b010000010010: io_out <= 8'b00000011;
		12'b010000010011: io_out <= 8'b01111101;
		12'b010000010100: io_out <= 8'b01011011;
		12'b010000010101: io_out <= 8'b10111000;
		12'b010000010110: io_out <= 8'b11110111;
		12'b010000010111: io_out <= 8'b11010100;
		12'b010000011000: io_out <= 8'b00010111;
		12'b010000011001: io_out <= 8'b01101101;
		12'b010000011010: io_out <= 8'b00011111;
		12'b010000011011: io_out <= 8'b10001010;
		12'b010000011100: io_out <= 8'b10110110;
		12'b010000011101: io_out <= 8'b00010110;
		12'b010000011110: io_out <= 8'b00111100;
		12'b010000011111: io_out <= 8'b00000011;
		12'b010000100000: io_out <= 8'b01100001;
		12'b010000100001: io_out <= 8'b01110110;
		12'b010000100010: io_out <= 8'b00000100;
		12'b010000100011: io_out <= 8'b01010110;
		12'b010000100100: io_out <= 8'b01111010;
		12'b010000100101: io_out <= 8'b10000001;
		12'b010000100110: io_out <= 8'b10000010;
		12'b010000100111: io_out <= 8'b00000011;
		12'b010000101000: io_out <= 8'b00111101;
		12'b010000101001: io_out <= 8'b10000100;
		12'b010000101010: io_out <= 8'b00101010;
		12'b010000101011: io_out <= 8'b10000111;
		12'b010000101100: io_out <= 8'b00110100;
		12'b010000101101: io_out <= 8'b00010010;
		12'b010000101110: io_out <= 8'b10001011;
		12'b010000101111: io_out <= 8'b00111110;
		12'b010000110000: io_out <= 8'b10001011;
		12'b010000110001: io_out <= 8'b10000011;
		12'b010000110010: io_out <= 8'b01000110;
		12'b010000110011: io_out <= 8'b01000110;
		12'b010000110100: io_out <= 8'b10001110;
		12'b010000110101: io_out <= 8'b00011101;
		12'b010000110110: io_out <= 8'b01011101;
		12'b010000110111: io_out <= 8'b00010001;
		12'b010000111000: io_out <= 8'b00111101;
		12'b010000111001: io_out <= 8'b00000001;
		12'b010000111010: io_out <= 8'b00000010;
		12'b010000111011: io_out <= 8'b01101101;
		12'b010000111100: io_out <= 8'b00111111;
		12'b010000111101: io_out <= 8'b00000010;
		12'b010000111110: io_out <= 8'b00000001;
		12'b010000111111: io_out <= 8'b10100010;
		12'b010001000000: io_out <= 8'b10100010;
		12'b010001000001: io_out <= 8'b10011110;
		12'b010001000010: io_out <= 8'b00100000;
		12'b010001000011: io_out <= 8'b00011101;
		12'b010001000100: io_out <= 8'b00100000;
		12'b010001000101: io_out <= 8'b10011100;
		12'b010001000110: io_out <= 8'b10100100;
		12'b010001000111: io_out <= 8'b01101000;
		12'b010001001000: io_out <= 8'b00000110;
		12'b010001001001: io_out <= 8'b10100001;
		12'b010001001010: io_out <= 8'b10100011;
		12'b010001001011: io_out <= 8'b10011101;
		12'b010001001100: io_out <= 8'b10001101;
		12'b010001001101: io_out <= 8'b01001010;
		12'b010001001110: io_out <= 8'b10100111;
		12'b010001001111: io_out <= 8'b10101001;
		12'b010001010000: io_out <= 8'b10100011;
		12'b010001010001: io_out <= 8'b00111101;
		12'b010001010010: io_out <= 8'b10010010;
		12'b010001010011: io_out <= 8'b10101110;
		12'b010001010100: io_out <= 8'b10110100;
		12'b010001010101: io_out <= 8'b01010011;
		12'b010001010110: io_out <= 8'b10110010;
		12'b010001010111: io_out <= 8'b10110111;
		12'b010001011000: io_out <= 8'b10100100;
		12'b010001011001: io_out <= 8'b01000110;
		12'b010001011010: io_out <= 8'b10111011;
		12'b010001011011: io_out <= 8'b10011101;
		12'b010001011100: io_out <= 8'b10000101;
		12'b010001011101: io_out <= 8'b00000100;
		12'b010001011110: io_out <= 8'b10101101;
		12'b010001011111: io_out <= 8'b10110111;
		12'b010001100000: io_out <= 8'b10010110;
		12'b010001100001: io_out <= 8'b10110011;
		12'b010001100010: io_out <= 8'b10100100;
		12'b010001100011: io_out <= 8'b11000000;
		12'b010001100100: io_out <= 8'b11000010;
		12'b010001100101: io_out <= 8'b10101110;
		12'b010001100110: io_out <= 8'b10010110;
		12'b010001100111: io_out <= 8'b00111100;
		12'b010001101000: io_out <= 8'b11001001;
		12'b010001101001: io_out <= 8'b11000111;
		12'b010001101010: io_out <= 8'b10111110;
		12'b010001101011: io_out <= 8'b11001010;
		12'b010001101100: io_out <= 8'b10001011;
		12'b010001101101: io_out <= 8'b11001100;
		12'b010001101110: io_out <= 8'b10000101;
		12'b010001101111: io_out <= 8'b11001000;
		12'b010001110000: io_out <= 8'b11001001;
		12'b010001110001: io_out <= 8'b10110101;
		12'b010001110010: io_out <= 8'b11010000;
		12'b010001110011: io_out <= 8'b10111000;
		12'b010001110100: io_out <= 8'b11010010;
		12'b010001110101: io_out <= 8'b10111110;
		12'b010001110110: io_out <= 8'b10011101;
		12'b010001110111: io_out <= 8'b10100001;
		12'b010001111000: io_out <= 8'b00111110;
		12'b010001111001: io_out <= 8'b11001000;
		12'b010001111010: io_out <= 8'b10100101;
		12'b010001111011: io_out <= 8'b10110001;
		12'b010001111100: io_out <= 8'b10110010;
		12'b010001111101: io_out <= 8'b11010011;
		12'b010001111110: io_out <= 8'b10111100;
		12'b010001111111: io_out <= 8'b11100010;
		12'b010010000000: io_out <= 8'b11010001;
		12'b010010000001: io_out <= 8'b00010111;
		12'b010010000010: io_out <= 8'b00011100;
		12'b010010000011: io_out <= 8'b00110000;
		12'b010010000100: io_out <= 8'b11000101;
		12'b010010000101: io_out <= 8'b11100011;
		12'b010010000110: io_out <= 8'b11001110;
		12'b010010000111: io_out <= 8'b01110110;
		12'b010010001000: io_out <= 8'b01001111;
		12'b010010001001: io_out <= 8'b11100001;
		12'b010010001010: io_out <= 8'b11101000;
		12'b010010001011: io_out <= 8'b11100100;
		12'b010010001100: io_out <= 8'b00101010;
		12'b010010001101: io_out <= 8'b11101100;
		12'b010010001110: io_out <= 8'b10111011;
		12'b010010001111: io_out <= 8'b11101110;
		12'b010010010000: io_out <= 8'b11000110;
		12'b010010010001: io_out <= 8'b11101011;
		12'b010010010010: io_out <= 8'b11001011;
		12'b010010010011: io_out <= 8'b11000011;
		12'b010010010100: io_out <= 8'b11010011;
		12'b010010010101: io_out <= 8'b10010111;
		12'b010010010110: io_out <= 8'b11000111;
		12'b010010010111: io_out <= 8'b11100001;
		12'b010010011000: io_out <= 8'b10011101;
		12'b010010011001: io_out <= 8'b10111011;
		12'b010010011010: io_out <= 8'b01111100;
		12'b010010011011: io_out <= 8'b11010010;
		12'b010010011100: io_out <= 8'b11111011;
		12'b010010011101: io_out <= 8'b11101000;
		12'b010010011110: io_out <= 8'b11111100;
		12'b010010011111: io_out <= 8'b01001001;
		12'b010010100000: io_out <= 8'b01001000;
		12'b010010100011: io_out <= 8'b00100001;
		12'b010010100100: io_out <= 8'b11111001;
		12'b010010100101: io_out <= 8'b00000100;
		12'b010010100110: io_out <= 8'b00000101;
		12'b010010100111: io_out <= 8'b00001101;
		12'b010010101011: io_out <= 8'b00101100;
		12'b010010110000: io_out <= 8'b00100000;
		12'b010010110010: io_out <= 8'b00100000;
		12'b010010110100: io_out <= 8'b10000010;
		12'b010010111000: io_out <= 8'b00110000;
		12'b010010111001: io_out <= 8'b00101010;
		12'b010010111010: io_out <= 8'b00011101;
		12'b010010111011: io_out <= 8'b01011111;
		12'b010010111100: io_out <= 8'b01001010;
		12'b010010111101: io_out <= 8'b01000010;
		12'b010010111110: io_out <= 8'b10010110;
		12'b010010111111: io_out <= 8'b01101000;
		12'b010011000000: io_out <= 8'b01100110;
		12'b010011000001: io_out <= 8'b10011111;
		12'b010011000010: io_out <= 8'b10011010;
		12'b010011000011: io_out <= 8'b10101001;
		12'b010011000100: io_out <= 8'b10101010;
		12'b010011000101: io_out <= 8'b10110001;
		12'b010011000110: io_out <= 8'b11001110;
		12'b010011000111: io_out <= 8'b10111011;
		12'b010011001000: io_out <= 8'b11000000;
		12'b010011001001: io_out <= 8'b11011110;
		12'b010011001010: io_out <= 8'b10000011;
		12'b010011001011: io_out <= 8'b01111100;
		12'b010011001100: io_out <= 8'b10000011;
		12'b010011001101: io_out <= 8'b00000011;
		12'b010011001110: io_out <= 8'b11011110;
		12'b010011001111: io_out <= 8'b01011000;
		12'b010011010000: io_out <= 8'b01100101;
		12'b010011010001: io_out <= 8'b11011010;
		12'b010011010011: io_out <= 8'b10000101;
		12'b010011010100: io_out <= 8'b11001000;
		12'b010011010101: io_out <= 8'b11011001;
		12'b010011010110: io_out <= 8'b00100010;
		12'b010011010111: io_out <= 8'b10110001;
		12'b010011011000: io_out <= 8'b10110010;
		12'b010011011001: io_out <= 8'b10101010;
		12'b010011011010: io_out <= 8'b01010111;
		12'b010011011011: io_out <= 8'b00011110;
		12'b010011011100: io_out <= 8'b11000111;
		12'b010011011101: io_out <= 8'b01011001;
		12'b010011011110: io_out <= 8'b00110101;
		12'b010011011111: io_out <= 8'b10001101;
		12'b010011100000: io_out <= 8'b10011011;
		12'b010011100001: io_out <= 8'b11000111;
		12'b010011100010: io_out <= 8'b00110001;
		12'b010011100011: io_out <= 8'b01100010;
		12'b010011100100: io_out <= 8'b10100100;
		12'b010011100101: io_out <= 8'b10000100;
		12'b010011100110: io_out <= 8'b00100000;
		12'b010011100111: io_out <= 8'b11011001;
		12'b010011101000: io_out <= 8'b01000001;
		12'b010011101001: io_out <= 8'b00100101;
		12'b010011101010: io_out <= 8'b10111100;
		12'b010011101011: io_out <= 8'b10101010;
		12'b010011101100: io_out <= 8'b10010110;
		12'b010011101101: io_out <= 8'b11010110;
		12'b010011101110: io_out <= 8'b01100110;
		12'b010011101111: io_out <= 8'b11011111;
		12'b010011110000: io_out <= 8'b00101011;
		12'b010011110001: io_out <= 8'b01011111;
		12'b010011110010: io_out <= 8'b00100011;
		12'b010011110011: io_out <= 8'b10110101;
		12'b010011110100: io_out <= 8'b11110110;
		12'b010011110101: io_out <= 8'b00010011;
		12'b010011110110: io_out <= 8'b00010011;
		12'b010011110111: io_out <= 8'b00001100;
		12'b010011111000: io_out <= 8'b10100101;
		12'b010011111001: io_out <= 8'b00100010;
		12'b010011111010: io_out <= 8'b00001100;
		12'b010011111011: io_out <= 8'b10001110;
		12'b010011111100: io_out <= 8'b10111110;
		12'b010011111101: io_out <= 8'b00011111;
		12'b010011111110: io_out <= 8'b11110000;
		12'b010011111111: io_out <= 8'b10010011;
		12'b010100000000: io_out <= 8'b11111011;
		12'b010100000001: io_out <= 8'b00001101;
		12'b010100000010: io_out <= 8'b00000100;
		12'b010100000011: io_out <= 8'b01010000;
		12'b010100000100: io_out <= 8'b11000001;
		12'b010100000101: io_out <= 8'b10000000;
		12'b010100000110: io_out <= 8'b10100111;
		12'b010100000111: io_out <= 8'b11101100;
		12'b010100001000: io_out <= 8'b00110001;
		12'b010100001001: io_out <= 8'b01110010;
		12'b010100001010: io_out <= 8'b00001100;
		12'b010100001011: io_out <= 8'b10000110;
		12'b010100001100: io_out <= 8'b11100100;
		12'b010100001101: io_out <= 8'b00011001;
		12'b010100001110: io_out <= 8'b00010101;
		12'b010100010000: io_out <= 8'b00101001;
		12'b010100010001: io_out <= 8'b11001001;
		12'b010100010010: io_out <= 8'b10001010;
		12'b010100010011: io_out <= 8'b11000111;
		12'b010100010100: io_out <= 8'b01110010;
		12'b010100010101: io_out <= 8'b00101100;
		12'b010100010110: io_out <= 8'b01111011;
		12'b010100010111: io_out <= 8'b10111111;
		12'b010100011000: io_out <= 8'b10010111;
		12'b010100011001: io_out <= 8'b10011001;
		12'b010100011010: io_out <= 8'b11001101;
		12'b010100011011: io_out <= 8'b11000000;
		12'b010100011100: io_out <= 8'b00100110;
		12'b010100011101: io_out <= 8'b10010111;
		12'b010100011110: io_out <= 8'b10011111;
		12'b010100011111: io_out <= 8'b11101000;
		12'b010100100000: io_out <= 8'b11010000;
		12'b010100100001: io_out <= 8'b11100101;
		12'b010100100010: io_out <= 8'b00101010;
		12'b010100100011: io_out <= 8'b01101011;
		12'b010100100100: io_out <= 8'b00011000;
		12'b010100100101: io_out <= 8'b11011111;
		12'b010100100110: io_out <= 8'b11110000;
		12'b010100100111: io_out <= 8'b01111000;
		12'b010100101000: io_out <= 8'b11001101;
		12'b010100101001: io_out <= 8'b10111110;
		12'b010100101010: io_out <= 8'b11011111;
		12'b010100101011: io_out <= 8'b11100010;
		12'b010100101100: io_out <= 8'b10100111;
		12'b010100101101: io_out <= 8'b01110001;
		12'b010100101110: io_out <= 8'b00101100;
		12'b010100101111: io_out <= 8'b01010101;
		12'b010100110000: io_out <= 8'b01001110;
		12'b010100110001: io_out <= 8'b01111000;
		12'b010100110010: io_out <= 8'b10000001;
		12'b010100110011: io_out <= 8'b00100100;
		12'b010100110100: io_out <= 8'b10000111;
		12'b010100110101: io_out <= 8'b00011001;
		12'b010100110110: io_out <= 8'b01111110;
		12'b010100110111: io_out <= 8'b01000111;
		12'b010100111000: io_out <= 8'b01100111;
		12'b010100111001: io_out <= 8'b10000110;
		12'b010100111010: io_out <= 8'b01000000;
		12'b010100111011: io_out <= 8'b01010101;
		12'b010100111100: io_out <= 8'b10001010;
		12'b010100111101: io_out <= 8'b01111001;
		12'b010100111110: io_out <= 8'b10001101;
		12'b010100111111: io_out <= 8'b01101001;
		12'b010101000000: io_out <= 8'b01110010;
		12'b010101000001: io_out <= 8'b00011000;
		12'b010101000010: io_out <= 8'b01111000;
		12'b010101000011: io_out <= 8'b10001100;
		12'b010101000100: io_out <= 8'b10001101;
		12'b010101000101: io_out <= 8'b10001111;
		12'b010101000110: io_out <= 8'b01000110;
		12'b010101000111: io_out <= 8'b01010001;
		12'b010101001000: io_out <= 8'b10010110;
		12'b010101001001: io_out <= 8'b10010111;
		12'b010101001010: io_out <= 8'b10010010;
		12'b010101001011: io_out <= 8'b01011011;
		12'b010101001100: io_out <= 8'b01010001;
		12'b010101001101: io_out <= 8'b00000001;
		12'b010101001110: io_out <= 8'b01011110;
		12'b010101001111: io_out <= 8'b01100101;
		12'b010101010000: io_out <= 8'b00000100;
		12'b010101010001: io_out <= 8'b01011101;
		12'b010101010010: io_out <= 8'b10011110;
		12'b010101010011: io_out <= 8'b00010010;
		12'b010101010100: io_out <= 8'b01010000;
		12'b010101010101: io_out <= 8'b00000001;
		12'b010101010110: io_out <= 8'b10101001;
		12'b010101010111: io_out <= 8'b10100001;
		12'b010101011000: io_out <= 8'b01011011;
		12'b010101011001: io_out <= 8'b00000100;
		12'b010101011010: io_out <= 8'b00000111;
		12'b010101011011: io_out <= 8'b00000010;
		12'b010101011100: io_out <= 8'b10101010;
		12'b010101011101: io_out <= 8'b01010000;
		12'b010101011110: io_out <= 8'b10011110;
		12'b010101011111: io_out <= 8'b10101111;
		12'b010101100000: io_out <= 8'b10101010;
		12'b010101100001: io_out <= 8'b10101001;
		12'b010101100010: io_out <= 8'b01010000;
		12'b010101100011: io_out <= 8'b01010011;
		12'b010101100100: io_out <= 8'b10101000;
		12'b010101100101: io_out <= 8'b10110100;
		12'b010101100110: io_out <= 8'b10011101;
		12'b010101100111: io_out <= 8'b01011111;
		12'b010101101000: io_out <= 8'b10110011;
		12'b010101101001: io_out <= 8'b10110100;
		12'b010101101010: io_out <= 8'b10100001;
		12'b010101101011: io_out <= 8'b01011101;
		12'b010101101100: io_out <= 8'b10111101;
		12'b010101101101: io_out <= 8'b10101011;
		12'b010101101110: io_out <= 8'b10000110;
		12'b010101101111: io_out <= 8'b10111100;
		12'b010101110000: io_out <= 8'b10111101;
		12'b010101110001: io_out <= 8'b10111111;
		12'b010101110010: io_out <= 8'b11000100;
		12'b010101110011: io_out <= 8'b10001101;
		12'b010101110100: io_out <= 8'b11000011;
		12'b010101110101: io_out <= 8'b10110000;
		12'b010101110110: io_out <= 8'b11000101;
		12'b010101110111: io_out <= 8'b10111001;
		12'b010101111000: io_out <= 8'b11000111;
		12'b010101111001: io_out <= 8'b11000000;
		12'b010101111010: io_out <= 8'b01010010;
		12'b010101111011: io_out <= 8'b10001011;
		12'b010101111100: io_out <= 8'b11001000;
		12'b010101111101: io_out <= 8'b11000001;
		12'b010101111110: io_out <= 8'b10000001;
		12'b010101111111: io_out <= 8'b11010000;
		12'b010110000000: io_out <= 8'b11001110;
		12'b010110000001: io_out <= 8'b01011100;
		12'b010110000010: io_out <= 8'b11001101;
		12'b010110000011: io_out <= 8'b10000110;
		12'b010110000100: io_out <= 8'b00000111;
		12'b010110000101: io_out <= 8'b11000000;
		12'b010110000110: io_out <= 8'b10100001;
		12'b010110000111: io_out <= 8'b01011100;
		12'b010110001000: io_out <= 8'b10111000;
		12'b010110001001: io_out <= 8'b11001011;
		12'b010110001010: io_out <= 8'b11010010;
		12'b010110001011: io_out <= 8'b11011001;
		12'b010110001100: io_out <= 8'b10101000;
		12'b010110001101: io_out <= 8'b10100000;
		12'b010110001110: io_out <= 8'b11000110;
		12'b010110001111: io_out <= 8'b01000110;
		12'b010110010000: io_out <= 8'b01101000;
		12'b010110010001: io_out <= 8'b11010000;
		12'b010110010010: io_out <= 8'b10111001;
		12'b010110010011: io_out <= 8'b11011100;
		12'b010110010100: io_out <= 8'b10111001;
		12'b010110010101: io_out <= 8'b10100011;
		12'b010110010110: io_out <= 8'b01000000;
		12'b010110010111: io_out <= 8'b11100101;
		12'b010110011000: io_out <= 8'b11100110;
		12'b010110011001: io_out <= 8'b11011111;
		12'b010110011010: io_out <= 8'b11101001;
		12'b010110011011: io_out <= 8'b00111101;
		12'b010110011100: io_out <= 8'b11101011;
		12'b010110011101: io_out <= 8'b11001001;
		12'b010110011110: io_out <= 8'b11011111;
		12'b010110011111: io_out <= 8'b11001110;
		12'b010110100000: io_out <= 8'b01011111;
		12'b010110100001: io_out <= 8'b10101110;
		12'b010110100010: io_out <= 8'b11011001;
		12'b010110100011: io_out <= 8'b11110001;
		12'b010110100100: io_out <= 8'b11110010;
		12'b010110100101: io_out <= 8'b10000000;
		12'b010110100110: io_out <= 8'b11101010;
		12'b010110100111: io_out <= 8'b10110110;
		12'b010110101000: io_out <= 8'b11010011;
		12'b010110101001: io_out <= 8'b11110000;
		12'b010110101010: io_out <= 8'b10110001;
		12'b010110101011: io_out <= 8'b00010011;
		12'b010110101100: io_out <= 8'b00001001;
		12'b010110101110: io_out <= 8'b00100001;
		12'b010110101111: io_out <= 8'b11111001;
		12'b010110110000: io_out <= 8'b00000100;
		12'b010110110001: io_out <= 8'b00000101;
		12'b010110110010: io_out <= 8'b00001101;
		12'b010110110110: io_out <= 8'b00101100;
		12'b010110111011: io_out <= 8'b00100000;
		12'b010110111101: io_out <= 8'b00100000;
		12'b010110111111: io_out <= 8'b10000010;
		12'b010111000011: io_out <= 8'b00110010;
		12'b010111000100: io_out <= 8'b00101100;
		12'b010111000101: io_out <= 8'b00100000;
		12'b010111000110: io_out <= 8'b01011101;
		12'b010111000111: io_out <= 8'b01001100;
		12'b010111001000: io_out <= 8'b01000101;
		12'b010111001001: io_out <= 8'b10011000;
		12'b010111001010: io_out <= 8'b01100111;
		12'b010111001011: io_out <= 8'b01100010;
		12'b010111001100: io_out <= 8'b10011101;
		12'b010111001101: io_out <= 8'b10011001;
		12'b010111001110: io_out <= 8'b10101000;
		12'b010111001111: io_out <= 8'b10101101;
		12'b010111010000: io_out <= 8'b10110100;
		12'b010111010001: io_out <= 8'b11010010;
		12'b010111010010: io_out <= 8'b10111011;
		12'b010111010011: io_out <= 8'b11000000;
		12'b010111010100: io_out <= 8'b11011111;
		12'b010111010101: io_out <= 8'b10010000;
		12'b010111010110: io_out <= 8'b01111110;
		12'b010111010111: io_out <= 8'b10000010;
		12'b010111011000: io_out <= 8'b00000011;
		12'b010111011001: io_out <= 8'b11111011;
		12'b010111011010: io_out <= 8'b00001000;
		12'b010111011011: io_out <= 8'b01100101;
		12'b010111011100: io_out <= 8'b10100101;
		12'b010111011101: io_out <= 8'b01101011;
		12'b010111011110: io_out <= 8'b10001100;
		12'b010111011111: io_out <= 8'b11001000;
		12'b010111100000: io_out <= 8'b01011001;
		12'b010111100001: io_out <= 8'b01101010;
		12'b010111100010: io_out <= 8'b10010001;
		12'b010111100011: io_out <= 8'b01110111;
		12'b010111100100: io_out <= 8'b10010010;
		12'b010111100101: io_out <= 8'b01101010;
		12'b010111100110: io_out <= 8'b00010100;
		12'b010111100111: io_out <= 8'b01010000;
		12'b010111101000: io_out <= 8'b00010000;
		12'b010111101001: io_out <= 8'b11010100;
		12'b010111101010: io_out <= 8'b01101000;
		12'b010111101011: io_out <= 8'b10011000;
		12'b010111101100: io_out <= 8'b01000101;
		12'b010111101101: io_out <= 8'b01001010;
		12'b010111101110: io_out <= 8'b01100000;
		12'b010111101111: io_out <= 8'b11110111;
		12'b010111110000: io_out <= 8'b10000001;
		12'b010111110001: io_out <= 8'b10010101;
		12'b010111110010: io_out <= 8'b01110011;
		12'b010111110011: io_out <= 8'b01101110;
		12'b010111110100: io_out <= 8'b01010111;
		12'b010111110101: io_out <= 8'b01000110;
		12'b010111110110: io_out <= 8'b00000010;
		12'b010111110111: io_out <= 8'b10010000;
		12'b010111111000: io_out <= 8'b11010111;
		12'b010111111001: io_out <= 8'b01111100;
		12'b010111111010: io_out <= 8'b11001101;
		12'b010111111011: io_out <= 8'b00100010;
		12'b010111111100: io_out <= 8'b00001101;
		12'b010111111101: io_out <= 8'b01111100;
		12'b010111111110: io_out <= 8'b00001001;
		12'b010111111111: io_out <= 8'b10111111;
		12'b011000000000: io_out <= 8'b00011011;
		12'b011000000001: io_out <= 8'b10011100;
		12'b011000000010: io_out <= 8'b10000111;
		12'b011000000011: io_out <= 8'b00010110;
		12'b011000000100: io_out <= 8'b00100001;
		12'b011000000101: io_out <= 8'b00001100;
		12'b011000000110: io_out <= 8'b00000100;
		12'b011000000111: io_out <= 8'b11001000;
		12'b011000001000: io_out <= 8'b00000001;
		12'b011000001001: io_out <= 8'b11000101;
		12'b011000001010: io_out <= 8'b11110100;
		12'b011000001011: io_out <= 8'b01011010;
		12'b011000001100: io_out <= 8'b11100001;
		12'b011000001101: io_out <= 8'b00010110;
		12'b011000001110: io_out <= 8'b00010101;
		12'b011000001111: io_out <= 8'b00100011;
		12'b011000010000: io_out <= 8'b01110010;
		12'b011000010001: io_out <= 8'b10101010;
		12'b011000010010: io_out <= 8'b10000100;
		12'b011000010011: io_out <= 8'b01000101;
		12'b011000010100: io_out <= 8'b00110101;
		12'b011000010101: io_out <= 8'b10011001;
		12'b011000010110: io_out <= 8'b11100111;
		12'b011000010111: io_out <= 8'b01010011;
		12'b011000011000: io_out <= 8'b00100111;
		12'b011000011001: io_out <= 8'b11100000;
		12'b011000011010: io_out <= 8'b01111001;
		12'b011000011011: io_out <= 8'b10101011;
		12'b011000011100: io_out <= 8'b10111110;
		12'b011000011101: io_out <= 8'b00010111;
		12'b011000011110: io_out <= 8'b01000011;
		12'b011000011111: io_out <= 8'b00101000;
		12'b011000100000: io_out <= 8'b00110010;
		12'b011000100001: io_out <= 8'b00010000;
		12'b011000100010: io_out <= 8'b10111010;
		12'b011000100011: io_out <= 8'b11011111;
		12'b011000100100: io_out <= 8'b10010011;
		12'b011000100101: io_out <= 8'b01101100;
		12'b011000100110: io_out <= 8'b00110011;
		12'b011000100111: io_out <= 8'b01110001;
		12'b011000101000: io_out <= 8'b00110110;
		12'b011000101001: io_out <= 8'b11001010;
		12'b011000101010: io_out <= 8'b11000110;
		12'b011000101011: io_out <= 8'b00101111;
		12'b011000101100: io_out <= 8'b00011000;
		12'b011000101101: io_out <= 8'b00011000;
		12'b011000101110: io_out <= 8'b00100011;
		12'b011000101111: io_out <= 8'b10101100;
		12'b011000110000: io_out <= 8'b01101110;
		12'b011000110001: io_out <= 8'b00001111;
		12'b011000110010: io_out <= 8'b10110011;
		12'b011000110011: io_out <= 8'b01111100;
		12'b011000110100: io_out <= 8'b10001110;
		12'b011000110101: io_out <= 8'b00100001;
		12'b011000110110: io_out <= 8'b01000101;
		12'b011000110111: io_out <= 8'b00111001;
		12'b011000111000: io_out <= 8'b01000010;
		12'b011000111001: io_out <= 8'b00100110;
		12'b011000111010: io_out <= 8'b01111011;
		12'b011000111011: io_out <= 8'b01111101;
		12'b011000111100: io_out <= 8'b01101010;
		12'b011000111101: io_out <= 8'b01101100;
		12'b011000111110: io_out <= 8'b01010110;
		12'b011000111111: io_out <= 8'b00010111;
		12'b011001000001: io_out <= 8'b00101000;
		12'b011001000010: io_out <= 8'b00011001;
		12'b011001000011: io_out <= 8'b01110010;
		12'b011001000100: io_out <= 8'b01000000;
		12'b011001000101: io_out <= 8'b01101010;
		12'b011001000110: io_out <= 8'b00010110;
		12'b011001000111: io_out <= 8'b10001001;
		12'b011001001000: io_out <= 8'b01101101;
		12'b011001001001: io_out <= 8'b10001011;
		12'b011001001010: io_out <= 8'b01101001;
		12'b011001001011: io_out <= 8'b01011000;
		12'b011001001100: io_out <= 8'b10001101;
		12'b011001001101: io_out <= 8'b10010000;
		12'b011001001110: io_out <= 8'b10000100;
		12'b011001001111: io_out <= 8'b01101100;
		12'b011001010000: io_out <= 8'b01110010;
		12'b011001010001: io_out <= 8'b00000010;
		12'b011001010010: io_out <= 8'b10001101;
		12'b011001010011: io_out <= 8'b10011011;
		12'b011001010100: io_out <= 8'b01010111;
		12'b011001010101: io_out <= 8'b00000100;
		12'b011001010110: io_out <= 8'b00000111;
		12'b011001010111: io_out <= 8'b01001001;
		12'b011001011000: io_out <= 8'b01011110;
		12'b011001011001: io_out <= 8'b01010011;
		12'b011001011010: io_out <= 8'b10011010;
		12'b011001011011: io_out <= 8'b10011011;
		12'b011001011100: io_out <= 8'b01110110;
		12'b011001011101: io_out <= 8'b10010000;
		12'b011001011110: io_out <= 8'b00110010;
		12'b011001011111: io_out <= 8'b01001000;
		12'b011001100000: io_out <= 8'b00000001;
		12'b011001100001: io_out <= 8'b01101000;
		12'b011001100010: io_out <= 8'b00111100;
		12'b011001100011: io_out <= 8'b01010011;
		12'b011001100100: io_out <= 8'b10101001;
		12'b011001100101: io_out <= 8'b10100011;
		12'b011001100110: io_out <= 8'b01000000;
		12'b011001100111: io_out <= 8'b00011111;
		12'b011001101000: io_out <= 8'b00011010;
		12'b011001101001: io_out <= 8'b10101000;
		12'b011001101010: io_out <= 8'b00000001;
		12'b011001101011: io_out <= 8'b10110011;
		12'b011001101100: io_out <= 8'b01001010;
		12'b011001101101: io_out <= 8'b10100001;
		12'b011001101110: io_out <= 8'b10110011;
		12'b011001101111: io_out <= 8'b10110011;
		12'b011001110000: io_out <= 8'b10101110;
		12'b011001110001: io_out <= 8'b10100100;
		12'b011001110010: io_out <= 8'b10110010;
		12'b011001110011: io_out <= 8'b10110111;
		12'b011001110100: io_out <= 8'b10011010;
		12'b011001110101: io_out <= 8'b01010101;
		12'b011001110110: io_out <= 8'b10111011;
		12'b011001110111: io_out <= 8'b10111001;
		12'b011001111000: io_out <= 8'b01110100;
		12'b011001111001: io_out <= 8'b10111011;
		12'b011001111010: io_out <= 8'b10110111;
		12'b011001111011: io_out <= 8'b10101101;
		12'b011001111100: io_out <= 8'b01000111;
		12'b011001111101: io_out <= 8'b00000010;
		12'b011001111110: io_out <= 8'b11000011;
		12'b011001111111: io_out <= 8'b11000000;
		12'b011010000000: io_out <= 8'b01000000;
		12'b011010000001: io_out <= 8'b11000110;
		12'b011010000010: io_out <= 8'b11000011;
		12'b011010000011: io_out <= 8'b10111100;
		12'b011010000100: io_out <= 8'b10100010;
		12'b011010000101: io_out <= 8'b11000111;
		12'b011010000110: io_out <= 8'b10100100;
		12'b011010000111: io_out <= 8'b00010010;
		12'b011010001000: io_out <= 8'b11001010;
		12'b011010001001: io_out <= 8'b11001011;
		12'b011010001010: io_out <= 8'b10101101;
		12'b011010001011: io_out <= 8'b11000010;
		12'b011010001100: io_out <= 8'b10101001;
		12'b011010001101: io_out <= 8'b00101111;
		12'b011010001110: io_out <= 8'b01101011;
		12'b011010001111: io_out <= 8'b01100111;
		12'b011010010000: io_out <= 8'b11010010;
		12'b011010010001: io_out <= 8'b10111000;
		12'b011010010010: io_out <= 8'b10101100;
		12'b011010010011: io_out <= 8'b11001011;
		12'b011010010100: io_out <= 8'b01111100;
		12'b011010010101: io_out <= 8'b00101111;
		12'b011010010110: io_out <= 8'b11010001;
		12'b011010010111: io_out <= 8'b11010010;
		12'b011010011000: io_out <= 8'b10100010;
		12'b011010011001: io_out <= 8'b11011111;
		12'b011010011010: io_out <= 8'b11001000;
		12'b011010011011: io_out <= 8'b00100111;
		12'b011010011100: io_out <= 8'b11011111;
		12'b011010011101: io_out <= 8'b11001011;
		12'b011010011110: io_out <= 8'b10100010;
		12'b011010011111: io_out <= 8'b01000111;
		12'b011010100000: io_out <= 8'b10111100;
		12'b011010100001: io_out <= 8'b10111010;
		12'b011010100010: io_out <= 8'b11011001;
		12'b011010100011: io_out <= 8'b11001100;
		12'b011010100100: io_out <= 8'b10100000;
		12'b011010100101: io_out <= 8'b11001010;
		12'b011010100110: io_out <= 8'b11100011;
		12'b011010100111: io_out <= 8'b10110001;
		12'b011010101000: io_out <= 8'b11101011;
		12'b011010101001: io_out <= 8'b11011010;
		12'b011010101010: io_out <= 8'b11101101;
		12'b011010101011: io_out <= 8'b10111000;
		12'b011010101100: io_out <= 8'b11101010;
		12'b011010101101: io_out <= 8'b11010011;
		12'b011010101110: io_out <= 8'b11100110;
		12'b011010101111: io_out <= 8'b10101000;
		12'b011010110000: io_out <= 8'b11011011;
		12'b011010110001: io_out <= 8'b11101111;
		12'b011010110010: io_out <= 8'b00010011;
		12'b011010110011: io_out <= 8'b11000110;
		12'b011010110100: io_out <= 8'b01101000;
		12'b011010110101: io_out <= 8'b11100101;
		12'b011010110110: io_out <= 8'b11111001;
		12'b011010110111: io_out <= 8'b10111000;
		12'b011010111000: io_out <= 8'b11011101;
		12'b011010111001: io_out <= 8'b01001000;
		12'b011010111010: io_out <= 8'b11110000;
		12'b011010111011: io_out <= 8'b10110011;
		12'b011010111100: io_out <= 8'b11000101;
		12'b011010111101: io_out <= 8'b11101110;
		12'b011010111110: io_out <= 8'b10011000;
		12'b011010111111: io_out <= 8'b10111110;
		12'b011011000000: io_out <= 8'b01111101;
		12'b011011000010: io_out <= 8'b00000111;
		12'b011011000011: io_out <= 8'b10000000;
		12'b011011000100: io_out <= 8'b10001011;
		12'b011011000101: io_out <= 8'b10000110;
		12'b011011000110: io_out <= 8'b11100100;
		12'b011011000111: io_out <= 8'b00011001;
		12'b011011001000: io_out <= 8'b00110100;
		12'b011011001001: io_out <= 8'b01101101;
		12'b011011001010: io_out <= 8'b00001011;
		12'b011011001011: io_out <= 8'b01110001;
		12'b011011001100: io_out <= 8'b00011101;
		12'b011011001101: io_out <= 8'b01110000;
		12'b011011001110: io_out <= 8'b10001000;
		12'b011011001111: io_out <= 8'b00110000;
		12'b011011010000: io_out <= 8'b01011011;
		12'b011011010001: io_out <= 8'b10111110;
		12'b011011010010: io_out <= 8'b01100111;
		12'b011011010011: io_out <= 8'b00001001;
		12'b011011010110: io_out <= 8'b00100001;
		12'b011011010111: io_out <= 8'b11111001;
		12'b011011011000: io_out <= 8'b00000100;
		12'b011011011001: io_out <= 8'b00000101;
		12'b011011011010: io_out <= 8'b00001101;
		12'b011011011110: io_out <= 8'b00101100;
		12'b011011100011: io_out <= 8'b00100000;
		12'b011011100101: io_out <= 8'b00100000;
		12'b011011100111: io_out <= 8'b10000010;
		12'b011011101011: io_out <= 8'b00110000;
		12'b011011101100: io_out <= 8'b00101010;
		12'b011011101101: io_out <= 8'b00011100;
		12'b011011101110: io_out <= 8'b01011100;
		12'b011011101111: io_out <= 8'b01001001;
		12'b011011110000: io_out <= 8'b01000010;
		12'b011011110001: io_out <= 8'b10010001;
		12'b011011110010: io_out <= 8'b01100001;
		12'b011011110011: io_out <= 8'b01011010;
		12'b011011110100: io_out <= 8'b10011100;
		12'b011011110101: io_out <= 8'b10010111;
		12'b011011110110: io_out <= 8'b10100111;
		12'b011011110111: io_out <= 8'b10101110;
		12'b011011111000: io_out <= 8'b10110101;
		12'b011011111001: io_out <= 8'b11010010;
		12'b011011111010: io_out <= 8'b10001101;
		12'b011011111011: io_out <= 8'b01111101;
		12'b011011111100: io_out <= 8'b10000010;
		12'b011100000000: io_out <= 8'b00000011;
		12'b011100000001: io_out <= 8'b11011100;
		12'b011100000010: io_out <= 8'b00001000;
		12'b011100000011: io_out <= 8'b10111010;
		12'b011100000100: io_out <= 8'b01011010;
		12'b011100000101: io_out <= 8'b01001110;
		12'b011100000110: io_out <= 8'b01100100;
		12'b011100000111: io_out <= 8'b01001000;
		12'b011100001000: io_out <= 8'b11101000;
		12'b011100001001: io_out <= 8'b00001010;
		12'b011100001010: io_out <= 8'b10111100;
		12'b011100001011: io_out <= 8'b10110111;
		12'b011100001100: io_out <= 8'b10110010;
		12'b011100001101: io_out <= 8'b01010101;
		12'b011100001110: io_out <= 8'b01010100;
		12'b011100001111: io_out <= 8'b10010100;
		12'b011100010000: io_out <= 8'b00100000;
		12'b011100010001: io_out <= 8'b01010001;
		12'b011100010010: io_out <= 8'b01100001;
		12'b011100010011: io_out <= 8'b00010111;
		12'b011100010100: io_out <= 8'b10110111;
		12'b011100010101: io_out <= 8'b00110001;
		12'b011100010110: io_out <= 8'b11010000;
		12'b011100010111: io_out <= 8'b00100000;
		12'b011100011000: io_out <= 8'b10101100;
		12'b011100011001: io_out <= 8'b11101011;
		12'b011100011010: io_out <= 8'b11110000;
		12'b011100011011: io_out <= 8'b10010000;
		12'b011100011100: io_out <= 8'b10011001;
		12'b011100011101: io_out <= 8'b11010110;
		12'b011100011110: io_out <= 8'b00111000;
		12'b011100011111: io_out <= 8'b10011110;
		12'b011100100000: io_out <= 8'b00101010;
		12'b011100100001: io_out <= 8'b10000000;
		12'b011100100010: io_out <= 8'b10000011;
		12'b011100100011: io_out <= 8'b01101000;
		12'b011100100100: io_out <= 8'b10111101;
		12'b011100100101: io_out <= 8'b00110000;
		12'b011100100110: io_out <= 8'b10111101;
		12'b011100100111: io_out <= 8'b00111101;
		12'b011100101000: io_out <= 8'b10110110;
		12'b011100101001: io_out <= 8'b00001001;
		12'b011100101010: io_out <= 8'b10100110;
		12'b011100101011: io_out <= 8'b01100010;
		12'b011100101100: io_out <= 8'b10000001;
		12'b011100101101: io_out <= 8'b10001001;
		12'b011100101110: io_out <= 8'b01001110;
		12'b011100101111: io_out <= 8'b11000000;
		12'b011100110000: io_out <= 8'b01010110;
		12'b011100110001: io_out <= 8'b10001000;
		12'b011100110010: io_out <= 8'b00110010;
		12'b011100110011: io_out <= 8'b00110010;
		12'b011100110100: io_out <= 8'b11111010;
		12'b011100110101: io_out <= 8'b01100110;
		12'b011100110110: io_out <= 8'b00010110;
		12'b011100110111: io_out <= 8'b11011100;
		12'b011100111000: io_out <= 8'b00110010;
		12'b011100111001: io_out <= 8'b01100110;
		12'b011100111010: io_out <= 8'b00100100;
		12'b011100111011: io_out <= 8'b10011100;
		12'b011100111100: io_out <= 8'b00010110;
		12'b011100111101: io_out <= 8'b00011111;
		12'b011100111110: io_out <= 8'b01101001;
		12'b011100111111: io_out <= 8'b00110101;
		12'b011101000000: io_out <= 8'b00010011;
		12'b011101000001: io_out <= 8'b11110011;
		12'b011101000010: io_out <= 8'b00010001;
		12'b011101000011: io_out <= 8'b00001101;
		12'b011101000100: io_out <= 8'b11010010;
		12'b011101000101: io_out <= 8'b11011100;
		12'b011101000110: io_out <= 8'b01010110;
		12'b011101000111: io_out <= 8'b01000100;
		12'b011101001000: io_out <= 8'b10010110;
		12'b011101001001: io_out <= 8'b00000001;
		12'b011101001010: io_out <= 8'b01110100;
		12'b011101001011: io_out <= 8'b01010001;
		12'b011101001100: io_out <= 8'b11101101;
		12'b011101001101: io_out <= 8'b01011000;
		12'b011101001110: io_out <= 8'b01100111;
		12'b011101001111: io_out <= 8'b11011101;
		12'b011101010000: io_out <= 8'b01100000;
		12'b011101010001: io_out <= 8'b11000010;
		12'b011101010010: io_out <= 8'b01101011;
		12'b011101010011: io_out <= 8'b00001010;
		12'b011101010100: io_out <= 8'b10010011;
		12'b011101010101: io_out <= 8'b01000111;
		12'b011101010110: io_out <= 8'b00010000;
		12'b011101010111: io_out <= 8'b00000100;
		12'b011101011000: io_out <= 8'b01101110;
		12'b011101011001: io_out <= 8'b11101010;
		12'b011101011010: io_out <= 8'b00111000;
		12'b011101011011: io_out <= 8'b11110001;
		12'b011101011100: io_out <= 8'b11000010;
		12'b011101011101: io_out <= 8'b10111010;
		12'b011101011110: io_out <= 8'b01001011;
		12'b011101011111: io_out <= 8'b01011001;
		12'b011101100000: io_out <= 8'b00000010;
		12'b011101100001: io_out <= 8'b01110010;
		12'b011101100010: io_out <= 8'b01010101;
		12'b011101100011: io_out <= 8'b01000101;
		12'b011101100100: io_out <= 8'b01110101;
		12'b011101100101: io_out <= 8'b00101011;
		12'b011101100110: io_out <= 8'b00000001;
		12'b011101100111: io_out <= 8'b10000111;
		12'b011101101000: io_out <= 8'b10000001;
		12'b011101101001: io_out <= 8'b00100001;
		12'b011101101010: io_out <= 8'b10000000;
		12'b011101101011: io_out <= 8'b10000001;
		12'b011101101100: io_out <= 8'b01110001;
		12'b011101101101: io_out <= 8'b10000101;
		12'b011101101110: io_out <= 8'b10000111;
		12'b011101101111: io_out <= 8'b10001111;
		12'b011101110000: io_out <= 8'b00110111;
		12'b011101110001: io_out <= 8'b00010001;
		12'b011101110010: io_out <= 8'b10000101;
		12'b011101110011: io_out <= 8'b10000000;
		12'b011101110100: io_out <= 8'b10001101;
		12'b011101110101: io_out <= 8'b01110101;
		12'b011101110110: io_out <= 8'b10001111;
		12'b011101110111: io_out <= 8'b10010111;
		12'b011101111000: io_out <= 8'b10001011;
		12'b011101111001: io_out <= 8'b01111101;
		12'b011101111010: io_out <= 8'b00000010;
		12'b011101111011: io_out <= 8'b00000110;
		12'b011101111100: io_out <= 8'b01110001;
		12'b011101111101: io_out <= 8'b00000110;
		12'b011101111110: io_out <= 8'b10010111;
		12'b011101111111: io_out <= 8'b10011111;
		12'b011110000000: io_out <= 8'b10011001;
		12'b011110000001: io_out <= 8'b10001111;
		12'b011110000010: io_out <= 8'b01100010;
		12'b011110000011: io_out <= 8'b01100011;
		12'b011110000100: io_out <= 8'b01110110;
		12'b011110000101: io_out <= 8'b10011111;
		12'b011110000110: io_out <= 8'b10010000;
		12'b011110000111: io_out <= 8'b10100001;
		12'b011110001000: io_out <= 8'b00000001;
		12'b011110001001: io_out <= 8'b10100011;
		12'b011110001010: io_out <= 8'b01011011;
		12'b011110001011: io_out <= 8'b10100101;
		12'b011110001100: io_out <= 8'b10100110;
		12'b011110001101: io_out <= 8'b01110111;
		12'b011110001110: io_out <= 8'b10001011;
		12'b011110001111: io_out <= 8'b10100010;
		12'b011110010000: io_out <= 8'b01110001;
		12'b011110010001: io_out <= 8'b10101100;
		12'b011110010010: io_out <= 8'b10100110;
		12'b011110010011: io_out <= 8'b10011010;
		12'b011110010100: io_out <= 8'b10101100;
		12'b011110010101: io_out <= 8'b10101010;
		12'b011110010110: io_out <= 8'b01000110;
		12'b011110010111: io_out <= 8'b10110010;
		12'b011110011000: io_out <= 8'b10101101;
		12'b011110011001: io_out <= 8'b10000110;
		12'b011110011010: io_out <= 8'b10000110;
		12'b011110011011: io_out <= 8'b10001000;
		12'b011110011100: io_out <= 8'b10000011;
		12'b011110011101: io_out <= 8'b00010000;
		12'b011110011110: io_out <= 8'b10111000;
		12'b011110011111: io_out <= 8'b10110011;
		12'b011110100000: io_out <= 8'b10000000;
		12'b011110100001: io_out <= 8'b10010000;
		12'b011110100010: io_out <= 8'b01101011;
		12'b011110100011: io_out <= 8'b10111111;
		12'b011110100100: io_out <= 8'b10011000;
		12'b011110100101: io_out <= 8'b11000001;
		12'b011110100110: io_out <= 8'b10010000;
		12'b011110100111: io_out <= 8'b10110110;
		12'b011110101000: io_out <= 8'b00100100;
		12'b011110101001: io_out <= 8'b11000100;
		12'b011110101010: io_out <= 8'b10001000;
		12'b011110101011: io_out <= 8'b00110111;
		12'b011110101100: io_out <= 8'b01111101;
		12'b011110101101: io_out <= 8'b10011000;
		12'b011110101110: io_out <= 8'b01000010;
		12'b011110101111: io_out <= 8'b00110000;
		12'b011110110000: io_out <= 8'b11001010;
		12'b011110110001: io_out <= 8'b01111110;
		12'b011110110010: io_out <= 8'b00010010;
		12'b011110110011: io_out <= 8'b01110111;
		12'b011110110100: io_out <= 8'b10100000;
		12'b011110110101: io_out <= 8'b11001111;
		12'b011110110110: io_out <= 8'b11001001;
		12'b011110110111: io_out <= 8'b10101101;
		12'b011110111000: io_out <= 8'b11001011;
		12'b011110111001: io_out <= 8'b10111010;
		12'b011110111010: io_out <= 8'b11010101;
		12'b011110111011: io_out <= 8'b11001000;
		12'b011110111100: io_out <= 8'b01111100;
		12'b011110111101: io_out <= 8'b11011000;
		12'b011110111110: io_out <= 8'b10101110;
		12'b011110111111: io_out <= 8'b01110110;
		12'b011111000000: io_out <= 8'b10100101;
		12'b011111000001: io_out <= 8'b10101100;
		12'b011111000010: io_out <= 8'b10011011;
		12'b011111000011: io_out <= 8'b01011011;
		12'b011111000100: io_out <= 8'b00000110;
		12'b011111000101: io_out <= 8'b10111011;
		12'b011111000110: io_out <= 8'b11011110;
		12'b011111000111: io_out <= 8'b10110000;
		12'b011111001000: io_out <= 8'b00010010;
		12'b011111001001: io_out <= 8'b10011100;
		12'b011111001010: io_out <= 8'b01101011;
		12'b011111001011: io_out <= 8'b00000011;
		12'b011111001100: io_out <= 8'b11100111;
		12'b011111001101: io_out <= 8'b11010100;
		12'b011111001110: io_out <= 8'b10101001;
		12'b011111001111: io_out <= 8'b10010101;
		12'b011111010000: io_out <= 8'b10111110;
		12'b011111010001: io_out <= 8'b11101101;
		12'b011111010010: io_out <= 8'b11100001;
		12'b011111010011: io_out <= 8'b11110000;
		12'b011111010100: io_out <= 8'b10010110;
		12'b011111010101: io_out <= 8'b11011000;
		12'b011111010110: io_out <= 8'b11100000;
		12'b011111010111: io_out <= 8'b10111100;
		12'b011111011000: io_out <= 8'b11110000;
		12'b011111011001: io_out <= 8'b11010001;
		12'b011111011010: io_out <= 8'b11110111;
		12'b011111011011: io_out <= 8'b01110111;
		12'b011111011100: io_out <= 8'b01110001;
		12'b011111011101: io_out <= 8'b00001001;
		12'b011111011111: io_out <= 8'b00100001;
		12'b011111100000: io_out <= 8'b11111001;
		12'b011111100001: io_out <= 8'b00000100;
		12'b011111100010: io_out <= 8'b00000101;
		12'b011111100011: io_out <= 8'b00011010;
		12'b011111100111: io_out <= 8'b00101100;
		12'b011111101100: io_out <= 8'b00100000;
		12'b011111101110: io_out <= 8'b00100000;
		12'b011111110000: io_out <= 8'b10000010;
		12'b011111110100: io_out <= 8'b00101111;
		12'b011111110101: io_out <= 8'b00101010;
		12'b011111110110: io_out <= 8'b00011100;
		12'b011111110111: io_out <= 8'b01011011;
		12'b011111111000: io_out <= 8'b01001000;
		12'b011111111001: io_out <= 8'b01000001;
		12'b011111111010: io_out <= 8'b10010101;
		12'b011111111011: io_out <= 8'b01100100;
		12'b011111111100: io_out <= 8'b01011101;
		12'b011111111101: io_out <= 8'b10011100;
		12'b011111111110: io_out <= 8'b10011000;
		12'b011111111111: io_out <= 8'b10101000;
		12'b100000000000: io_out <= 8'b10101001;
		12'b100000000001: io_out <= 8'b10110000;
		12'b100000000010: io_out <= 8'b11001110;
		12'b100000000011: io_out <= 8'b10111010;
		12'b100000000100: io_out <= 8'b11000000;
		12'b100000000101: io_out <= 8'b11011110;
		12'b100000000110: io_out <= 8'b10010111;
		12'b100000000111: io_out <= 8'b01111110;
		12'b100000001000: io_out <= 8'b10000010;
		12'b100000001001: io_out <= 8'b00000011;
		12'b100000001010: io_out <= 8'b11101010;
		12'b100000001011: io_out <= 8'b01011000;
		12'b100000001100: io_out <= 8'b01100101;
		12'b100000001101: io_out <= 8'b10101010;
		12'b100000001110: io_out <= 8'b11110000;
		12'b100000001111: io_out <= 8'b10000101;
		12'b100000010000: io_out <= 8'b11001000;
		12'b100000010001: io_out <= 8'b11011001;
		12'b100000010010: io_out <= 8'b00100010;
		12'b100000010011: io_out <= 8'b10110001;
		12'b100000010100: io_out <= 8'b10110010;
		12'b100000010101: io_out <= 8'b10110001;
		12'b100000010110: io_out <= 8'b00000010;
		12'b100000010111: io_out <= 8'b00011111;
		12'b100000011000: io_out <= 8'b10010100;
		12'b100000011001: io_out <= 8'b01000011;
		12'b100000011010: io_out <= 8'b00111000;
		12'b100000011011: io_out <= 8'b01011100;
		12'b100000011100: io_out <= 8'b01001101;
		12'b100000011101: io_out <= 8'b00110110;
		12'b100000011110: io_out <= 8'b10010001;
		12'b100000011111: io_out <= 8'b10011100;
		12'b100000100000: io_out <= 8'b00000111;
		12'b100000100001: io_out <= 8'b00101100;
		12'b100000100010: io_out <= 8'b00100101;
		12'b100000100011: io_out <= 8'b00110001;
		12'b100000100100: io_out <= 8'b00001000;
		12'b100000100101: io_out <= 8'b00110000;
		12'b100000100110: io_out <= 8'b01001100;
		12'b100000100111: io_out <= 8'b10011110;
		12'b100000101000: io_out <= 8'b10110100;
		12'b100000101001: io_out <= 8'b10110011;
		12'b100000101010: io_out <= 8'b11011010;
		12'b100000101011: io_out <= 8'b11100101;
		12'b100000101100: io_out <= 8'b00011011;
		12'b100000101101: io_out <= 8'b00001011;
		12'b100000101110: io_out <= 8'b10100011;
		12'b100000101111: io_out <= 8'b00110010;
		12'b100000110000: io_out <= 8'b11010011;
		12'b100000110001: io_out <= 8'b00011001;
		12'b100000110010: io_out <= 8'b10001000;
		12'b100000110011: io_out <= 8'b01101101;
		12'b100000110100: io_out <= 8'b01000101;
		12'b100000110101: io_out <= 8'b10001000;
		12'b100000110110: io_out <= 8'b10001001;
		12'b100000110111: io_out <= 8'b01100110;
		12'b100000111000: io_out <= 8'b00010101;
		12'b100000111001: io_out <= 8'b10100000;
		12'b100000111010: io_out <= 8'b01000100;
		12'b100000111011: io_out <= 8'b01110101;
		12'b100000111100: io_out <= 8'b00100011;
		12'b100000111101: io_out <= 8'b11000010;
		12'b100000111110: io_out <= 8'b01000100;
		12'b100000111111: io_out <= 8'b10000111;
		12'b100001000000: io_out <= 8'b01010011;
		12'b100001000001: io_out <= 8'b01010010;
		12'b100001000010: io_out <= 8'b10111010;
		12'b100001000011: io_out <= 8'b01101100;
		12'b100001000100: io_out <= 8'b11011110;
		12'b100001000101: io_out <= 8'b00100010;
		12'b100001000110: io_out <= 8'b01001111;
		12'b100001000111: io_out <= 8'b11010001;
		12'b100001001000: io_out <= 8'b11101000;
		12'b100001001001: io_out <= 8'b10010010;
		12'b100001001010: io_out <= 8'b11000001;
		12'b100001001011: io_out <= 8'b11010000;
		12'b100001001100: io_out <= 8'b00011000;
		12'b100001001101: io_out <= 8'b10011101;
		12'b100001001110: io_out <= 8'b01001111;
		12'b100001001111: io_out <= 8'b10001000;
		12'b100001010000: io_out <= 8'b01110111;
		12'b100001010001: io_out <= 8'b10101100;
		12'b100001010010: io_out <= 8'b01010001;
		12'b100001010011: io_out <= 8'b10111011;
		12'b100001010100: io_out <= 8'b00010101;
		12'b100001010101: io_out <= 8'b01010110;
		12'b100001010110: io_out <= 8'b01000001;
		12'b100001010111: io_out <= 8'b01011011;
		12'b100001011000: io_out <= 8'b11110110;
		12'b100001011001: io_out <= 8'b01001010;
		12'b100001011010: io_out <= 8'b01111101;
		12'b100001011011: io_out <= 8'b11101001;
		12'b100001011100: io_out <= 8'b11001000;
		12'b100001011101: io_out <= 8'b11000110;
		12'b100001011110: io_out <= 8'b10100101;
		12'b100001011111: io_out <= 8'b01010101;
		12'b100001100000: io_out <= 8'b01111010;
		12'b100001100001: io_out <= 8'b01001011;
		12'b100001100010: io_out <= 8'b01110001;
		12'b100001100011: io_out <= 8'b00011010;
		12'b100001100100: io_out <= 8'b11011011;
		12'b100001100101: io_out <= 8'b01111110;
		12'b100001100110: io_out <= 8'b01000111;
		12'b100001100111: io_out <= 8'b10111011;
		12'b100001101000: io_out <= 8'b11011001;
		12'b100001101001: io_out <= 8'b00100001;
		12'b100001101010: io_out <= 8'b01000000;
		12'b100001101011: io_out <= 8'b01101110;
		12'b100001101100: io_out <= 8'b00010100;
		12'b100001101101: io_out <= 8'b00101101;
		12'b100001101110: io_out <= 8'b00100000;
		12'b100001101111: io_out <= 8'b01000110;
		12'b100001110000: io_out <= 8'b01011010;
		12'b100001110001: io_out <= 8'b00000010;
		12'b100001110010: io_out <= 8'b01010001;
		12'b100001110011: io_out <= 8'b00010100;
		12'b100001110100: io_out <= 8'b01001010;
		12'b100001110101: io_out <= 8'b00100110;
		12'b100001110110: io_out <= 8'b00010011;
		12'b100001110111: io_out <= 8'b00111010;
		12'b100001111000: io_out <= 8'b00000001;
		12'b100001111001: io_out <= 8'b00000001;
		12'b100001111010: io_out <= 8'b01100100;
		12'b100001111011: io_out <= 8'b00100001;
		12'b100001111100: io_out <= 8'b00000111;
		12'b100001111101: io_out <= 8'b01000110;
		12'b100001111110: io_out <= 8'b10001100;
		12'b100001111111: io_out <= 8'b01001010;
		12'b100010000000: io_out <= 8'b10001111;
		12'b100010000001: io_out <= 8'b10010000;
		12'b100010000010: io_out <= 8'b10010001;
		12'b100010000011: io_out <= 8'b00000100;
		12'b100010000100: io_out <= 8'b00000111;
		12'b100010000101: io_out <= 8'b01011011;
		12'b100010000110: io_out <= 8'b00111011;
		12'b100010000111: io_out <= 8'b00000010;
		12'b100010001000: io_out <= 8'b10010110;
		12'b100010001001: io_out <= 8'b00110100;
		12'b100010001010: io_out <= 8'b00000010;
		12'b100010001011: io_out <= 8'b10011001;
		12'b100010001100: io_out <= 8'b10011001;
		12'b100010001101: io_out <= 8'b10001001;
		12'b100010001110: io_out <= 8'b10011100;
		12'b100010001111: io_out <= 8'b01000101;
		12'b100010010000: io_out <= 8'b00110001;
		12'b100010010001: io_out <= 8'b10011010;
		12'b100010010010: io_out <= 8'b10100000;
		12'b100010010011: io_out <= 8'b00010011;
		12'b100010010100: io_out <= 8'b10100011;
		12'b100010010101: io_out <= 8'b10100011;
		12'b100010010110: io_out <= 8'b10011110;
		12'b100010010111: io_out <= 8'b00110000;
		12'b100010011000: io_out <= 8'b10100100;
		12'b100010011001: io_out <= 8'b10101010;
		12'b100010011010: io_out <= 8'b01000101;
		12'b100010011011: io_out <= 8'b10101100;
		12'b100010011100: io_out <= 8'b10101101;
		12'b100010011101: io_out <= 8'b10011110;
		12'b100010011110: io_out <= 8'b10110000;
		12'b100010011111: io_out <= 8'b10101010;
		12'b100010100000: io_out <= 8'b10100010;
		12'b100010100001: io_out <= 8'b10110011;
		12'b100010100010: io_out <= 8'b10010000;
		12'b100010100011: io_out <= 8'b10101110;
		12'b100010100100: io_out <= 8'b10110110;
		12'b100010100101: io_out <= 8'b10100000;
		12'b100010100110: io_out <= 8'b10111000;
		12'b100010100111: io_out <= 8'b10111001;
		12'b100010101000: io_out <= 8'b10101000;
		12'b100010101001: io_out <= 8'b10101111;
		12'b100010101010: io_out <= 8'b10111010;
		12'b100010101011: io_out <= 8'b10101010;
		12'b100010101100: io_out <= 8'b00000011;
		12'b100010101101: io_out <= 8'b10111001;
		12'b100010101110: io_out <= 8'b10100100;
		12'b100010101111: io_out <= 8'b10101111;
		12'b100010110000: io_out <= 8'b11000001;
		12'b100010110001: io_out <= 8'b10101001;
		12'b100010110010: io_out <= 8'b10000010;
		12'b100010110011: io_out <= 8'b00010010;
		12'b100010110100: io_out <= 8'b10111110;
		12'b100010110101: io_out <= 8'b11000101;
		12'b100010110110: io_out <= 8'b11000111;
		12'b100010110111: io_out <= 8'b10101101;
		12'b100010111000: io_out <= 8'b10110111;
		12'b100010111001: io_out <= 8'b11000101;
		12'b100010111010: io_out <= 8'b11000110;
		12'b100010111011: io_out <= 8'b10010001;
		12'b100010111100: io_out <= 8'b11001111;
		12'b100010111101: io_out <= 8'b10111101;
		12'b100010111110: io_out <= 8'b11010001;
		12'b100010111111: io_out <= 8'b10100100;
		12'b100011000000: io_out <= 8'b11010011;
		12'b100011000001: io_out <= 8'b10111100;
		12'b100011000010: io_out <= 8'b10001100;
		12'b100011000011: io_out <= 8'b11001100;
		12'b100011000100: io_out <= 8'b10111111;
		12'b100011000101: io_out <= 8'b10100010;
		12'b100011000110: io_out <= 8'b11001100;
		12'b100011000111: io_out <= 8'b10011111;
		12'b100011001000: io_out <= 8'b10010110;
		12'b100011001001: io_out <= 8'b10010100;
		12'b100011001010: io_out <= 8'b11010001;
		12'b100011001011: io_out <= 8'b00111011;
		12'b100011001100: io_out <= 8'b11011000;
		12'b100011001101: io_out <= 8'b10111010;
		12'b100011001110: io_out <= 8'b10000001;
		12'b100011001111: io_out <= 8'b11011010;
		12'b100011010000: io_out <= 8'b11001101;
		12'b100011010001: io_out <= 8'b00101111;
		12'b100011010010: io_out <= 8'b00101111;
		12'b100011010011: io_out <= 8'b11100100;
		12'b100011010100: io_out <= 8'b10010001;
		12'b100011010101: io_out <= 8'b00111100;
		12'b100011010110: io_out <= 8'b11010101;
		12'b100011010111: io_out <= 8'b10110011;
		12'b100011011000: io_out <= 8'b10010010;
		12'b100011011001: io_out <= 8'b11011101;
		12'b100011011010: io_out <= 8'b10101100;
		12'b100011011011: io_out <= 8'b11101101;
		12'b100011011100: io_out <= 8'b10010110;
		12'b100011011101: io_out <= 8'b10011000;
		12'b100011011110: io_out <= 8'b11000110;
		12'b100011011111: io_out <= 8'b11101010;
		12'b100011100000: io_out <= 8'b11011000;
		12'b100011100001: io_out <= 8'b10111110;
		12'b100011100010: io_out <= 8'b11011111;
		12'b100011100011: io_out <= 8'b11010000;
		12'b100011100100: io_out <= 8'b11100010;
		12'b100011100101: io_out <= 8'b10111010;
		12'b100011100110: io_out <= 8'b10010100;
		12'b100011100111: io_out <= 8'b00110010;
		12'b100011101000: io_out <= 8'b10110001;
		12'b100011101001: io_out <= 8'b11011011;
		12'b100011101010: io_out <= 8'b01101000;
		12'b100011101011: io_out <= 8'b00001001;
		12'b100011101100: io_out <= 8'b10001011;
		12'b100011101101: io_out <= 8'b01110101;
		12'b100011101110: io_out <= 8'b00100010;
		12'b100011101111: io_out <= 8'b10100000;
		12'b100011110000: io_out <= 8'b00110100;
		12'b100011110001: io_out <= 8'b01001000;
		12'b100011110010: io_out <= 8'b10110001;
		12'b100011110011: io_out <= 8'b00010010;
		12'b100011110110: io_out <= 8'b00100001;
		12'b100011110111: io_out <= 8'b11111001;
		12'b100011111000: io_out <= 8'b00000100;
		12'b100011111001: io_out <= 8'b00000101;
		12'b100011111010: io_out <= 8'b00001101;
		12'b100011111110: io_out <= 8'b00101100;
		12'b100100000011: io_out <= 8'b00100000;
		12'b100100000101: io_out <= 8'b00100000;
		12'b100100000111: io_out <= 8'b10000010;
		12'b100100001011: io_out <= 8'b00110000;
		12'b100100001100: io_out <= 8'b00101011;
		12'b100100001101: io_out <= 8'b00011111;
		12'b100100001110: io_out <= 8'b01011001;
		12'b100100001111: io_out <= 8'b01001001;
		12'b100100010000: io_out <= 8'b01000010;
		12'b100100010001: io_out <= 8'b10011001;
		12'b100100010010: io_out <= 8'b01101000;
		12'b100100010011: io_out <= 8'b01100101;
		12'b100100010100: io_out <= 8'b10011111;
		12'b100100010101: io_out <= 8'b10011010;
		12'b100100010110: io_out <= 8'b10101001;
		12'b100100010111: io_out <= 8'b10101110;
		12'b100100011000: io_out <= 8'b10110100;
		12'b100100011001: io_out <= 8'b11010000;
		12'b100100011010: io_out <= 8'b10010101;
		12'b100100011011: io_out <= 8'b01111101;
		12'b100100011100: io_out <= 8'b10000011;
		12'b100100100000: io_out <= 8'b00000011;
		12'b100100100001: io_out <= 8'b11101010;
		12'b100100100010: io_out <= 8'b00001000;
		12'b100100100011: io_out <= 8'b10110101;
		12'b100100100100: io_out <= 8'b10111010;
		12'b100100100101: io_out <= 8'b10100101;
		12'b100100100110: io_out <= 8'b00100100;
		12'b100100100111: io_out <= 8'b01001010;
		12'b100100101000: io_out <= 8'b01010111;
		12'b100100101001: io_out <= 8'b10100100;
		12'b100100101010: io_out <= 8'b00100101;
		12'b100100101011: io_out <= 8'b01001100;
		12'b100100101100: io_out <= 8'b10000001;
		12'b100100101101: io_out <= 8'b01000110;
		12'b100100101110: io_out <= 8'b11101011;
		12'b100100101111: io_out <= 8'b11101101;
		12'b100100110000: io_out <= 8'b11010001;
		12'b100100110001: io_out <= 8'b00100110;
		12'b100100110010: io_out <= 8'b01100110;
		12'b100100110011: io_out <= 8'b10100011;
		12'b100100110100: io_out <= 8'b11010011;
		12'b100100110101: io_out <= 8'b01011100;
		12'b100100110110: io_out <= 8'b10010001;
		12'b100100110111: io_out <= 8'b10000011;
		12'b100100111000: io_out <= 8'b10100110;
		12'b100100111001: io_out <= 8'b10001111;
		12'b100100111010: io_out <= 8'b11010110;
		12'b100100111011: io_out <= 8'b01000010;
		12'b100100111100: io_out <= 8'b10001011;
		12'b100100111101: io_out <= 8'b11100101;
		12'b100100111110: io_out <= 8'b10000001;
		12'b100100111111: io_out <= 8'b01100010;
		12'b100101000000: io_out <= 8'b11011101;
		12'b100101000001: io_out <= 8'b00111110;
		12'b100101000010: io_out <= 8'b10101111;
		12'b100101000011: io_out <= 8'b00110111;
		12'b100101000100: io_out <= 8'b00001100;
		12'b100101000101: io_out <= 8'b11000010;
		12'b100101000110: io_out <= 8'b10001110;
		12'b100101000111: io_out <= 8'b01110101;
		12'b100101001000: io_out <= 8'b10011110;
		12'b100101001001: io_out <= 8'b01010000;
		12'b100101001010: io_out <= 8'b11001101;
		12'b100101001011: io_out <= 8'b10100110;
		12'b100101001100: io_out <= 8'b11100010;
		12'b100101001101: io_out <= 8'b00001001;
		12'b100101001110: io_out <= 8'b10001110;
		12'b100101001111: io_out <= 8'b10111101;
		12'b100101010000: io_out <= 8'b10001001;
		12'b100101010001: io_out <= 8'b10101010;
		12'b100101010010: io_out <= 8'b01000110;
		12'b100101010011: io_out <= 8'b00100000;
		12'b100101010100: io_out <= 8'b01101110;
		12'b100101010101: io_out <= 8'b10001010;
		12'b100101010110: io_out <= 8'b10111101;
		12'b100101010111: io_out <= 8'b01011101;
		12'b100101011000: io_out <= 8'b01010010;
		12'b100101011001: io_out <= 8'b01010110;
		12'b100101011010: io_out <= 8'b00011001;
		12'b100101011011: io_out <= 8'b10001110;
		12'b100101011100: io_out <= 8'b10011110;
		12'b100101011101: io_out <= 8'b00011100;
		12'b100101011110: io_out <= 8'b11000010;
		12'b100101011111: io_out <= 8'b01101110;
		12'b100101100000: io_out <= 8'b11101011;
		12'b100101100001: io_out <= 8'b01011011;
		12'b100101100010: io_out <= 8'b01001101;
		12'b100101100011: io_out <= 8'b10101100;
		12'b100101100100: io_out <= 8'b00001100;
		12'b100101100101: io_out <= 8'b10011100;
		12'b100101100110: io_out <= 8'b10010110;
		12'b100101100111: io_out <= 8'b11011011;
		12'b100101101000: io_out <= 8'b00001101;
		12'b100101101001: io_out <= 8'b01111110;
		12'b100101101010: io_out <= 8'b00110010;
		12'b100101101011: io_out <= 8'b00111000;
		12'b100101101101: io_out <= 8'b01101011;
		12'b100101101110: io_out <= 8'b11001100;
		12'b100101101111: io_out <= 8'b00110101;
		12'b100101110000: io_out <= 8'b10100000;
		12'b100101110001: io_out <= 8'b11001100;
		12'b100101110010: io_out <= 8'b10111111;
		12'b100101110011: io_out <= 8'b01011111;
		12'b100101110100: io_out <= 8'b00011000;
		12'b100101110101: io_out <= 8'b00010011;
		12'b100101110110: io_out <= 8'b00100001;
		12'b100101110111: io_out <= 8'b00001111;
		12'b100101111000: io_out <= 8'b11010110;
		12'b100101111001: io_out <= 8'b10101001;
		12'b100101111010: io_out <= 8'b00001111;
		12'b100101111011: io_out <= 8'b10001011;
		12'b100101111100: io_out <= 8'b10100100;
		12'b100101111101: io_out <= 8'b10101110;
		12'b100101111110: io_out <= 8'b01110011;
		12'b100101111111: io_out <= 8'b11011111;
		12'b100110000000: io_out <= 8'b00010110;
		12'b100110000001: io_out <= 8'b01001110;
		12'b100110000010: io_out <= 8'b01001100;
		12'b100110000011: io_out <= 8'b00010110;
		12'b100110000100: io_out <= 8'b01110110;
		12'b100110000101: io_out <= 8'b01101110;
		12'b100110000110: io_out <= 8'b00010011;
		12'b100110000111: io_out <= 8'b00101000;
		12'b100110001000: io_out <= 8'b01010110;
		12'b100110001001: io_out <= 8'b01111001;
		12'b100110001010: io_out <= 8'b10000100;
		12'b100110001011: io_out <= 8'b01011100;
		12'b100110001100: io_out <= 8'b01010011;
		12'b100110001101: io_out <= 8'b01011110;
		12'b100110001110: io_out <= 8'b10000001;
		12'b100110001111: io_out <= 8'b00011011;
		12'b100110010000: io_out <= 8'b10001010;
		12'b100110010001: io_out <= 8'b00010001;
		12'b100110010010: io_out <= 8'b00000110;
		12'b100110010011: io_out <= 8'b01100100;
		12'b100110010100: io_out <= 8'b01001000;
		12'b100110010101: io_out <= 8'b00000010;
		12'b100110010110: io_out <= 8'b10001110;
		12'b100110010111: io_out <= 8'b10001111;
		12'b100110011000: io_out <= 8'b00101000;
		12'b100110011001: io_out <= 8'b01000111;
		12'b100110011010: io_out <= 8'b01110110;
		12'b100110011011: io_out <= 8'b01000111;
		12'b100110011100: io_out <= 8'b00000001;
		12'b100110011101: io_out <= 8'b01001000;
		12'b100110011110: io_out <= 8'b10001111;
		12'b100110011111: io_out <= 8'b00100010;
		12'b100110100000: io_out <= 8'b00101011;
		12'b100110100001: io_out <= 8'b10011100;
		12'b100110100010: io_out <= 8'b10011101;
		12'b100110100011: io_out <= 8'b01011011;
		12'b100110100100: io_out <= 8'b00010001;
		12'b100110100101: io_out <= 8'b00000010;
		12'b100110100110: io_out <= 8'b00000001;
		12'b100110100111: io_out <= 8'b10100111;
		12'b100110101000: io_out <= 8'b10100011;
		12'b100110101001: io_out <= 8'b00010111;
		12'b100110101010: io_out <= 8'b01000011;
		12'b100110101011: io_out <= 8'b00010010;
		12'b100110101100: io_out <= 8'b00000110;
		12'b100110101101: io_out <= 8'b10100110;
		12'b100110101110: io_out <= 8'b10101000;
		12'b100110101111: io_out <= 8'b10010110;
		12'b100110110000: io_out <= 8'b10010011;
		12'b100110110001: io_out <= 8'b10100101;
		12'b100110110010: io_out <= 8'b10101000;
		12'b100110110011: io_out <= 8'b10100111;
		12'b100110110100: io_out <= 8'b10010110;
		12'b100110110101: io_out <= 8'b10010111;
		12'b100110110110: io_out <= 8'b10110010;
		12'b100110110111: io_out <= 8'b10110011;
		12'b100110111000: io_out <= 8'b10010101;
		12'b100110111001: io_out <= 8'b01001000;
		12'b100110111010: io_out <= 8'b10110011;
		12'b100110111011: io_out <= 8'b10011101;
		12'b100110111100: io_out <= 8'b10110110;
		12'b100110111101: io_out <= 8'b01011010;
		12'b100110111110: io_out <= 8'b10111011;
		12'b100110111111: io_out <= 8'b10110100;
		12'b100111000000: io_out <= 8'b10111001;
		12'b100111000001: io_out <= 8'b10111011;
		12'b100111000010: io_out <= 8'b10110101;
		12'b100111000011: io_out <= 8'b10010111;
		12'b100111000100: io_out <= 8'b10101110;
		12'b100111000101: io_out <= 8'b10111111;
		12'b100111000110: io_out <= 8'b10010101;
		12'b100111000111: io_out <= 8'b11000110;
		12'b100111001000: io_out <= 8'b10000000;
		12'b100111001001: io_out <= 8'b00010110;
		12'b100111001010: io_out <= 8'b11000101;
		12'b100111001011: io_out <= 8'b11000010;
		12'b100111001100: io_out <= 8'b11000111;
		12'b100111001101: io_out <= 8'b10111011;
		12'b100111001110: io_out <= 8'b10000110;
		12'b100111001111: io_out <= 8'b10001110;
		12'b100111010000: io_out <= 8'b11001011;
		12'b100111010001: io_out <= 8'b10111000;
		12'b100111010010: io_out <= 8'b10111001;
		12'b100111010011: io_out <= 8'b10100010;
		12'b100111010100: io_out <= 8'b10111100;
		12'b100111010101: io_out <= 8'b11000100;
		12'b100111010110: io_out <= 8'b10111111;
		12'b100111010111: io_out <= 8'b10101111;
		12'b100111011000: io_out <= 8'b01001000;
		12'b100111011001: io_out <= 8'b01011011;
		12'b100111011010: io_out <= 8'b10101110;
		12'b100111011011: io_out <= 8'b11000011;
		12'b100111011100: io_out <= 8'b01011110;
		12'b100111011101: io_out <= 8'b11010001;
		12'b100111011110: io_out <= 8'b11010010;
		12'b100111011111: io_out <= 8'b10011010;
		12'b100111100000: io_out <= 8'b01010010;
		12'b100111100001: io_out <= 8'b10110100;
		12'b100111100010: io_out <= 8'b10110110;
		12'b100111100011: io_out <= 8'b11011110;
		12'b100111100100: io_out <= 8'b11011000;
		12'b100111100101: io_out <= 8'b11011001;
		12'b100111100110: io_out <= 8'b00111100;
		12'b100111100111: io_out <= 8'b10101000;
		12'b100111101000: io_out <= 8'b01110111;
		12'b100111101001: io_out <= 8'b11010000;
		12'b100111101010: io_out <= 8'b11010111;
		12'b100111101011: io_out <= 8'b11011000;
		12'b100111101100: io_out <= 8'b11000000;
		12'b100111101101: io_out <= 8'b11011011;
		12'b100111101110: io_out <= 8'b11100011;
		12'b100111101111: io_out <= 8'b11100100;
		12'b100111110000: io_out <= 8'b11000000;
		12'b100111110001: io_out <= 8'b11000110;
		12'b100111110010: io_out <= 8'b11001111;
		12'b100111110011: io_out <= 8'b01011110;
		12'b100111110100: io_out <= 8'b10010011;
		12'b100111110101: io_out <= 8'b11100111;
		12'b100111110110: io_out <= 8'b11000110;
		12'b100111110111: io_out <= 8'b11010001;
		12'b100111111000: io_out <= 8'b01000111;
		12'b100111111001: io_out <= 8'b10111101;
		12'b100111111010: io_out <= 8'b11110101;
		12'b100111111011: io_out <= 8'b11100100;
		12'b100111111100: io_out <= 8'b11010100;
		12'b100111111101: io_out <= 8'b10001101;
		12'b100111111110: io_out <= 8'b10110110;
		12'b100111111111: io_out <= 8'b11011010;
		12'b101000000000: io_out <= 8'b11101011;
		12'b101000000001: io_out <= 8'b10001010;
		12'b101000000010: io_out <= 8'b01110001;
		12'b101000000011: io_out <= 8'b10110011;
		12'b101000000100: io_out <= 8'b10110101;
		12'b101000000101: io_out <= 8'b11101111;
		12'b101000000110: io_out <= 8'b10011010;
		12'b101000000111: io_out <= 8'b10101110;
		12'b101000001000: io_out <= 8'b01010011;
		12'b101000001001: io_out <= 8'b10110110;
		12'b101000001010: io_out <= 8'b00010010;
		12'b101000001101: io_out <= 8'b00100001;
		12'b101000001110: io_out <= 8'b11111001;
		12'b101000001111: io_out <= 8'b00000100;
		12'b101000010000: io_out <= 8'b00000101;
		12'b101000010001: io_out <= 8'b00001101;
		12'b101000010011: io_out <= 8'b00000111;
		12'b101000010101: io_out <= 8'b00101100;
		12'b101000011010: io_out <= 8'b00100000;
		12'b101000011100: io_out <= 8'b00100000;
		12'b101000011110: io_out <= 8'b10000010;
		12'b101000011111: io_out <= 8'b00110001;
		12'b101000100000: io_out <= 8'b00101100;
		12'b101000100001: io_out <= 8'b00100001;
		12'b101000100010: io_out <= 8'b01100101;
		12'b101000100011: io_out <= 8'b01010110;
		12'b101000100100: io_out <= 8'b01010011;
		12'b101000100101: io_out <= 8'b01010001;
		12'b101000100110: io_out <= 8'b00111110;
		12'b101000100111: io_out <= 8'b00110100;
		12'b101000101000: io_out <= 8'b10010101;
		12'b101000101001: io_out <= 8'b01100101;
		12'b101000101010: io_out <= 8'b01100000;
		12'b101000101011: io_out <= 8'b10011110;
		12'b101000101100: io_out <= 8'b10011010;
		12'b101000101101: io_out <= 8'b10101010;
		12'b101000101110: io_out <= 8'b10101100;
		12'b101000101111: io_out <= 8'b10110010;
		12'b101000110000: io_out <= 8'b11001111;
		12'b101000110001: io_out <= 8'b10111011;
		12'b101000110010: io_out <= 8'b11000000;
		12'b101000110011: io_out <= 8'b11011110;
		12'b101000110111: io_out <= 8'b00000011;
		12'b101000111000: io_out <= 8'b11100011;
		12'b101000111001: io_out <= 8'b01011000;
		12'b101000111010: io_out <= 8'b01100101;
		12'b101000111011: io_out <= 8'b10101010;
		12'b101000111100: io_out <= 8'b11000110;
		12'b101000111101: io_out <= 8'b10000101;
		12'b101000111110: io_out <= 8'b11001000;
		12'b101000111111: io_out <= 8'b11011001;
		12'b101001000000: io_out <= 8'b11100010;
		12'b101001000001: io_out <= 8'b10111100;
		12'b101001000010: io_out <= 8'b00101110;
		12'b101001000011: io_out <= 8'b10101111;
		12'b101001000100: io_out <= 8'b10100111;
		12'b101001000101: io_out <= 8'b00101110;
		12'b101001000110: io_out <= 8'b01101101;
		12'b101001000111: io_out <= 8'b10011110;
		12'b101001001000: io_out <= 8'b11100100;
		12'b101001001001: io_out <= 8'b01110000;
		12'b101001001010: io_out <= 8'b00001101;
		12'b101001001011: io_out <= 8'b00000100;
		12'b101001001100: io_out <= 8'b10000110;
		12'b101001001101: io_out <= 8'b00100111;
		12'b101001001110: io_out <= 8'b01101010;
		12'b101001001111: io_out <= 8'b00011100;
		12'b101001010000: io_out <= 8'b01000111;
		12'b101001010001: io_out <= 8'b11000011;
		12'b101001010010: io_out <= 8'b01110110;
		12'b101001010011: io_out <= 8'b10011101;
		12'b101001010100: io_out <= 8'b01101000;
		12'b101001010101: io_out <= 8'b11000001;
		12'b101001010110: io_out <= 8'b00010110;
		12'b101001010111: io_out <= 8'b11001010;
		12'b101001011000: io_out <= 8'b01100010;
		12'b101001011001: io_out <= 8'b10010101;
		12'b101001011010: io_out <= 8'b00011100;
		12'b101001011011: io_out <= 8'b00010011;
		12'b101001011100: io_out <= 8'b01111001;
		12'b101001011101: io_out <= 8'b01001000;
		12'b101001011110: io_out <= 8'b11011100;
		12'b101001011111: io_out <= 8'b10011111;
		12'b101001100000: io_out <= 8'b10011101;
		12'b101001100001: io_out <= 8'b01100100;
		12'b101001100010: io_out <= 8'b10000000;
		12'b101001100011: io_out <= 8'b00010011;
		12'b101001100100: io_out <= 8'b01011110;
		12'b101001100101: io_out <= 8'b01011110;
		12'b101001100110: io_out <= 8'b10111100;
		12'b101001100111: io_out <= 8'b01001010;
		12'b101001101000: io_out <= 8'b01101100;
		12'b101001101001: io_out <= 8'b00010000;
		12'b101001101010: io_out <= 8'b01101000;
		12'b101001101011: io_out <= 8'b00010010;
		12'b101001101100: io_out <= 8'b00111111;
		12'b101001101101: io_out <= 8'b00111110;
		12'b101001101110: io_out <= 8'b10000010;
		12'b101001101111: io_out <= 8'b10101001;
		12'b101001110000: io_out <= 8'b10110100;
		12'b101001110001: io_out <= 8'b10001000;
		12'b101001110010: io_out <= 8'b00110000;
		12'b101001110011: io_out <= 8'b10011011;
		12'b101001110100: io_out <= 8'b11001110;
		12'b101001110101: io_out <= 8'b00101000;
		12'b101001110110: io_out <= 8'b00101111;
		12'b101001110111: io_out <= 8'b01011000;
		12'b101001111000: io_out <= 8'b01100001;
		12'b101001111001: io_out <= 8'b00110000;
		12'b101001111010: io_out <= 8'b00001000;
		12'b101001111011: io_out <= 8'b10000011;
		12'b101001111100: io_out <= 8'b10110000;
		12'b101001111101: io_out <= 8'b00111000;
		12'b101001111110: io_out <= 8'b10100000;
		12'b101001111111: io_out <= 8'b10001101;
		12'b101010000000: io_out <= 8'b10011000;
		12'b101010000001: io_out <= 8'b10010101;
		12'b101010000010: io_out <= 8'b11001001;
		12'b101010000011: io_out <= 8'b10001110;
		12'b101010000100: io_out <= 8'b01111000;
		12'b101010000101: io_out <= 8'b10101101;
		12'b101010000110: io_out <= 8'b01001101;
		12'b101010000111: io_out <= 8'b00100110;
		12'b101010001000: io_out <= 8'b01001001;
		12'b101010001001: io_out <= 8'b11101001;
		12'b101010001010: io_out <= 8'b11100001;
		12'b101010001011: io_out <= 8'b00111010;
		12'b101010001100: io_out <= 8'b11011100;
		12'b101010001101: io_out <= 8'b10011110;
		12'b101010001110: io_out <= 8'b10100101;
		12'b101010001111: io_out <= 8'b01000010;
		12'b101010010000: io_out <= 8'b11110011;
		12'b101010010001: io_out <= 8'b01100111;
		12'b101010010010: io_out <= 8'b11111101;
		12'b101010010011: io_out <= 8'b10001110;
		12'b101010010100: io_out <= 8'b01100111;
		12'b101010010101: io_out <= 8'b01010011;
		12'b101010010110: io_out <= 8'b11001010;
		12'b101010010111: io_out <= 8'b01010000;
		12'b101010011000: io_out <= 8'b01111101;
		12'b101010011001: io_out <= 8'b01001100;
		12'b101010011010: io_out <= 8'b01111010;
		12'b101010011011: io_out <= 8'b01011011;
		12'b101010011100: io_out <= 8'b01101101;
		12'b101010011101: io_out <= 8'b00110010;
		12'b101010011110: io_out <= 8'b00111110;
		12'b101010011111: io_out <= 8'b01100011;
		12'b101010100000: io_out <= 8'b10000100;
		12'b101010100001: io_out <= 8'b10000110;
		12'b101010100010: io_out <= 8'b10001011;
		12'b101010100011: io_out <= 8'b01110011;
		12'b101010100100: io_out <= 8'b10001011;
		12'b101010100101: io_out <= 8'b10001110;
		12'b101010100110: io_out <= 8'b01111001;
		12'b101010100111: io_out <= 8'b01010111;
		12'b101010101000: io_out <= 8'b10001110;
		12'b101010101001: io_out <= 8'b01010001;
		12'b101010101010: io_out <= 8'b01001100;
		12'b101010101011: io_out <= 8'b00000010;
		12'b101010101100: io_out <= 8'b00000001;
		12'b101010101101: io_out <= 8'b01101100;
		12'b101010101110: io_out <= 8'b00000001;
		12'b101010110000: io_out <= 8'b10010101;
		12'b101010110001: io_out <= 8'b01100100;
		12'b101010110010: io_out <= 8'b10010010;
		12'b101010110011: io_out <= 8'b01100000;
		12'b101010110100: io_out <= 8'b00000001;
		12'b101010110101: io_out <= 8'b00000010;
		12'b101010111000: io_out <= 8'b01100100;
		12'b101010111001: io_out <= 8'b01100010;
		12'b101010111010: io_out <= 8'b00000100;
		12'b101010111011: io_out <= 8'b10011000;
		12'b101010111100: io_out <= 8'b10100000;
		12'b101010111101: io_out <= 8'b10011001;
		12'b101010111110: io_out <= 8'b10011011;
		12'b101010111111: io_out <= 8'b10001011;
		12'b101011000000: io_out <= 8'b10011111;
		12'b101011000001: io_out <= 8'b10100110;
		12'b101011000010: io_out <= 8'b10100010;
		12'b101011000011: io_out <= 8'b01100010;
		12'b101011000100: io_out <= 8'b10101010;
		12'b101011000101: io_out <= 8'b10100110;
		12'b101011000110: io_out <= 8'b10100001;
		12'b101011000111: io_out <= 8'b10001011;
		12'b101011001000: io_out <= 8'b10100101;
		12'b101011001001: io_out <= 8'b10101111;
		12'b101011001010: io_out <= 8'b10011010;
		12'b101011001011: io_out <= 8'b01001101;
		12'b101011001100: io_out <= 8'b10101111;
		12'b101011001101: io_out <= 8'b10101011;
		12'b101011001110: io_out <= 8'b00011000;
		12'b101011001111: io_out <= 8'b00111110;
		12'b101011010000: io_out <= 8'b10110010;
		12'b101011010001: io_out <= 8'b10100110;
		12'b101011010010: io_out <= 8'b10110100;
		12'b101011010011: io_out <= 8'b10111010;
		12'b101011010100: io_out <= 8'b10110111;
		12'b101011010101: io_out <= 8'b10000110;
		12'b101011010110: io_out <= 8'b10111101;
		12'b101011010111: io_out <= 8'b00000010;
		12'b101011011000: io_out <= 8'b10111100;
		12'b101011011001: io_out <= 8'b10110110;
		12'b101011011010: io_out <= 8'b10100000;
		12'b101011011011: io_out <= 8'b00000010;
		12'b101011011100: io_out <= 8'b10110001;
		12'b101011011101: io_out <= 8'b10111011;
		12'b101011011110: io_out <= 8'b10010110;
		12'b101011011111: io_out <= 8'b01011000;
		12'b101011100000: io_out <= 8'b10110101;
		12'b101011100001: io_out <= 8'b11000011;
		12'b101011100010: io_out <= 8'b10110000;
		12'b101011100011: io_out <= 8'b01101101;
		12'b101011100100: io_out <= 8'b10110010;
		12'b101011100101: io_out <= 8'b10010110;
		12'b101011100110: io_out <= 8'b01010111;
		12'b101011100111: io_out <= 8'b01011000;
		12'b101011101000: io_out <= 8'b11001011;
		12'b101011101001: io_out <= 8'b11001100;
		12'b101011101010: io_out <= 8'b01011010;
		12'b101011101011: io_out <= 8'b10110010;
		12'b101011101100: io_out <= 8'b01100011;
		12'b101011101101: io_out <= 8'b11001001;
		12'b101011101110: io_out <= 8'b11010010;
		12'b101011101111: io_out <= 8'b10101000;
		12'b101011110000: io_out <= 8'b01010001;
		12'b101011110001: io_out <= 8'b10101010;
		12'b101011110010: io_out <= 8'b00000010;
		12'b101011110011: io_out <= 8'b10101101;
		12'b101011110100: io_out <= 8'b10010101;
		12'b101011110101: io_out <= 8'b11000001;
		12'b101011110110: io_out <= 8'b11010010;
		12'b101011110111: io_out <= 8'b11000101;
		12'b101011111000: io_out <= 8'b11010100;
		12'b101011111001: io_out <= 8'b11011111;
		12'b101011111010: io_out <= 8'b11011110;
		12'b101011111011: io_out <= 8'b10101011;
		12'b101011111100: io_out <= 8'b11000001;
		12'b101011111101: io_out <= 8'b10101110;
		12'b101011111110: io_out <= 8'b10110110;
		12'b101011111111: io_out <= 8'b11011001;
		12'b101100000000: io_out <= 8'b00011110;
		12'b101100000001: io_out <= 8'b10111010;
		12'b101100000010: io_out <= 8'b11100111;
		12'b101100000011: io_out <= 8'b11100110;
		12'b101100000100: io_out <= 8'b11100111;
		12'b101100000101: io_out <= 8'b10101111;
		12'b101100000110: io_out <= 8'b11101001;
		12'b101100000111: io_out <= 8'b00010111;
		12'b101100001000: io_out <= 8'b10111101;
		12'b101100001001: io_out <= 8'b10110011;
		12'b101100001010: io_out <= 8'b10011110;
		12'b101100001011: io_out <= 8'b11101110;
		12'b101100001100: io_out <= 8'b10111110;
		12'b101100001101: io_out <= 8'b10001000;
		12'b101100001110: io_out <= 8'b11110101;
		12'b101100001111: io_out <= 8'b11000100;
		12'b101100010000: io_out <= 8'b01001101;
		12'b101100010001: io_out <= 8'b11111000;
		12'b101100010010: io_out <= 8'b11010011;
		12'b101100010011: io_out <= 8'b10111001;
		12'b101100010100: io_out <= 8'b11110100;
		12'b101100010101: io_out <= 8'b10110110;
		12'b101100010110: io_out <= 8'b10011010;
		12'b101100010111: io_out <= 8'b11111011;
		12'b101100011000: io_out <= 8'b10111000;
		12'b101100011001: io_out <= 8'b01001101;
		12'b101100011010: io_out <= 8'b01001000;
		12'b101100011101: io_out <= 8'b00111011;
		default: io_out <= 8'b00000000;
	endcase;
end

endmodule
